//bus_control_tb.v
//Author: RndMnkIII. 19/07/2021. (@RndMnkIII).
//---------------------------------------------------------
//iverilog -o bus_control_tb.vvp DFF2.v k053326_D21.v k053327_D20.v bus_control.v bus_control_tb.v
//vvp bus_control_tb.vvp -lxt2
//gtkwave bus_control_tb.lxt&
`default_nettype none
`timescale 1 ns/ 10 ps //time-unit = 1 ns, precision = 1 ps

module bus_control_tb;
    //SYSCLK=48Mhz, period 20.832ns; 12Mhz, period 83.333ns; 3Mhz period 333.33ns
	parameter TS = 10.416;
	parameter T64 = TS * 64;
	parameter TS56 = TS * 56;
	parameter TS40 = TS * 40;
	parameter TS33 = TS * 33;
	parameter TS32 = TS * 32;
	parameter TS29 = TS * 29;
	parameter TS23 = TS * 23;
	parameter TS20 = TS * 20;
	parameter TS17 = TS * 17;
	parameter TS16 = TS * 16;
	parameter TS14 = TS * 14;
	parameter TS13 = TS * 13;
	parameter TS11 = TS * 11;
	parameter TS10 = TS * 10;
	parameter TS8 = TS * 8;
	parameter TS5 = TS * 5;
	parameter TS4 = TS * 4;
	parameter TS3 = TS * 3;
	parameter TS2 = TS * 2;
	
	reg [16:0] x,y;

	reg AS, BK4, INIT;
	reg WOCO, RMRD;
	reg SYSCLK, CK12, CKE, CKQ;
	reg [15:0] ADDR;
	wire PROG, BANK, WORK, OBJCS, VRAMCS, CRAMCS, IOCS, DTAC, NCK12;
    
    reg NCLK12, RESETb;
    reg [7:0] DATA;
    reg RWb, AS2, DTAC2, VRAMCS2;
    
    reg tmp;
	always @(*) begin
        tmp = ~NCLK12;
        CK12 = tmp;
    end
    //CK12 = ~NCLK12; 
	BusControl ABC(.BK4(BK4), .INIT(INIT), .ADDR(ADDR), .WOCO(WOCO), .RMRD(RMRD), 
	                     .CE(CKE), .CQ(CKQ), .CLK12(CK12), .RWb(RWb),
						 .PROG(PROG), .BANK(BANK), .WORK(WORK), .OBJCS(OBJCS), .VRAMCS(VRAMCS), .CRAMCS(CRAMCS), .IOCS(IOCS), 
						 .AS(AS2), .DTAC(DTAC),
						 .CLK12n(NCK12));			 

	initial
	begin
		//INIT=1'b0;
		//#TS16
		INIT=1'b1;
		//RWb=1'b1;
	end
	
	
	//VRAMCS test
	// initial //RWb timing
	// begin
		// RWb=1'b1;
		// #TS4;
		// for (x=16'h4000; x <= 16'h7fff; x= x + 16'h0001)
		// begin
			
			// RWb=1'b1;
			// #TS8;
			// RWb=1'b0;
			// #TS23;
			// RWb=1'b1;
			// #TS;
		// end
	// end
	// initial //AS timing
	// begin
		// AS=1'b1;
		// #TS4;
		// for (x=16'h4000; x <= 16'h7fff; x= x + 16'h0001)
		// begin
			
			// AS=1'b1;
			// #TS10;
			// AS=1'b0;
			// #TS20;
			// AS=1'b1;
			// #TS2;
		// end
	// end
	
	// initial //ADDR timing
	// begin
		// ADDR = 16'hFFFF; 
		// #TS4;
		// for (y=16'h4000; y <= 16'h7fff; y= y + 16'h0001)
		// begin
			// ADDR = y[15:0];
			// #TS32;
		// end
	// end
	
	initial
	begin
		BK4 = 1'b0;
		RMRD = 1'b0;
		WOCO = 1'b0;
	end
	

	// always
	// begin
		// SYSCLK = 1'b0;
		// #TS; //high for 10.416 ns
		// SYSCLK = 1'b1;
		// #TS; //low for 10.416 ns
	// end

	// always
	// begin
		// //period 83.333ns
		// CK12 = 1'b0;
		// #TS2;
		// CK12 = 1'b1;
		// #TS2;
	// end
	
	// always
	// begin
		// CKE = 1'b0;
		// #TS8;
		// CKE = 1'b1;
		// #TS8;
	// end
	
	// always
	// begin
		// CKQ = 1'b0;
		// #TS4;
		// CKQ = 1'b1;
		// #TS8;
		// CKQ = 1'b0;
		// #TS4;
	// end
	
	initial
	begin
		$dumpfile ("bus_control_tb.lxt");
		$dumpvars (0, bus_control_tb); //0 all variables included
		//#46418500 $finish;
	end
    
    initial
begin
    NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #22.5; SYSCLK = 1'b0;
    #22.5; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b0;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; NCLK12 = 1'b1;
    SYSCLK = 1'b1;
    #20.0; SYSCLK = 1'b0;
    #20.0; 
end
initial
begin
    CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #170.0; CKE = 1'b0;
    #160.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;
    #160.0; CKE = 1'b0;
    #170.0; CKE = 1'b1;

end
initial
begin
    CKQ = 1'b0;
    #70.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #170.0; CKQ = 1'b0;
    #160.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;
    #170.0; CKQ = 1'b1;
    #160.0; CKQ = 1'b0;

end
initial
begin
    RESETb = 1'b1;

end
initial
begin
    ADDR = 16'h1EE2;
    #70.0; ADDR = 16'h1EE3;
    #400.0; ADDR = 16'h00AB;
    #10.0; ADDR = 16'h81AF;
    #400.0; ADDR = 16'h81A0;
    #10.0; ADDR = 16'h81B0;
    #650.0; ADDR = 16'h81A9;
    #410.0; ADDR = 16'h81AA;
    #410.0; ADDR = 16'h81AB;
    #400.0; ADDR = 16'h81A9;
    #10.0; ADDR = 16'h81AC;
    #400.0; ADDR = 16'h8880;
    #10.0; ADDR = 16'h1EC2;
    #490.0; ADDR = 16'h1EC3;
    #400.0; ADDR = 16'h04C3;
    #10.0; ADDR = 16'h81AD;
    #400.0; ADDR = 16'h81AC;
    #10.0; ADDR = 16'h81AE;
    #410.0; ADDR = 16'h81AF;
    #160.0; ADDR = 16'h1EE2;
    #580.0; ADDR = 16'h1EE3;
    #400.0; ADDR = 16'h81AF;
    #410.0; ADDR = 16'h81A0;
    #10.0; ADDR = 16'h81B0;
    #640.0; ADDR = 16'h81A0;
    #10.0; ADDR = 16'h81A9;
    #400.0; ADDR = 16'h81A8;
    #10.0; ADDR = 16'h81AA;
    #410.0; ADDR = 16'h81AB;
    #400.0; ADDR = 16'h81A8;
    #10.0; ADDR = 16'h81AC;
    #400.0; ADDR = 16'h1E80;
    #10.0; ADDR = 16'h1EC2;
    #490.0; ADDR = 16'h1EC3;
    #400.0; ADDR = 16'h01AD;
    #10.0; ADDR = 16'h81AD;
    #400.0; ADDR = 16'h81AC;
    #10.0; ADDR = 16'h81AE;
    #410.0; ADDR = 16'h81AF;
    #150.0; ADDR = 16'h1AA2;
    #10.0; ADDR = 16'h1EE2;
    #570.0; ADDR = 16'h1EE3;
    #400.0; ADDR = 16'h06E3;
    #10.0; ADDR = 16'h81AF;
    #400.0; ADDR = 16'h81A3;
    #10.0; ADDR = 16'h81B0;
    #650.0; ADDR = 16'h81A0;
    #10.0; ADDR = 16'h81A9;
    #400.0; ADDR = 16'h81A8;
    #10.0; ADDR = 16'h81AA;
    #400.0; ADDR = 16'h81AB;
    #410.0; ADDR = 16'h81AC;
    #400.0; ADDR = 16'h80AC;
    #10.0; ADDR = 16'h1EC2;
    #490.0; ADDR = 16'h1EC3;
    #400.0; ADDR = 16'h16C3;
    #10.0; ADDR = 16'h81AD;
    #410.0; ADDR = 16'h81AE;
    #410.0; ADDR = 16'h81AF;
    #160.0; ADDR = 16'h1EA2;
    #10.0; ADDR = 16'h1EE2;
    #570.0; ADDR = 16'h1EE3;
    #400.0; ADDR = 16'h01AF;
    #10.0; ADDR = 16'h81AF;
    #400.0; ADDR = 16'h81A0;
    #10.0; ADDR = 16'h81B0;
    #650.0; ADDR = 16'h81A9;
    #410.0; ADDR = 16'h81AA;
    #410.0; ADDR = 16'h81AB;
    #400.0; ADDR = 16'h81A8;
    #10.0; ADDR = 16'h81AC;
    #400.0; ADDR = 16'h1880;
    #10.0; ADDR = 16'h1EC2;
    #490.0; ADDR = 16'h1EC3;
    #400.0; ADDR = 16'h00C3;
    #10.0; ADDR = 16'h81AD;
    #400.0; ADDR = 16'h81AC;
    #10.0; ADDR = 16'h81AE;
    #410.0; ADDR = 16'h81AF;
    #160.0; ADDR = 16'h1EE2;
    #570.0; ADDR = 16'h1EE3;
    #410.0; ADDR = 16'h81AF;
    #410.0; ADDR = 16'h81A0;
    #10.0; ADDR = 16'h81B0;
    #640.0; ADDR = 16'h81A0;
    #10.0; ADDR = 16'h81A9;
    #400.0; ADDR = 16'h81A8;
    #10.0; ADDR = 16'h81AA;
    #410.0; ADDR = 16'h81AB;
    #400.0; ADDR = 16'h81A8;
    #10.0; ADDR = 16'h81AC;
    #400.0; ADDR = 16'h1E80;
    #10.0; ADDR = 16'h1EC2;
    #490.0; ADDR = 16'h1EC3;
    #400.0; ADDR = 16'h01AD;
    #10.0; ADDR = 16'h81AD;
    #400.0; ADDR = 16'h81AC;
    #10.0; ADDR = 16'h81AE;
    #410.0; ADDR = 16'h81AF;
    #150.0; ADDR = 16'h18A2;
    #10.0; ADDR = 16'h1EE2;
    #570.0; ADDR = 16'h1EE3;
    #400.0; ADDR = 16'h06E3;
    #10.0; ADDR = 16'h81AF;
    #410.0; ADDR = 16'h81B0;
    #650.0; ADDR = 16'h81A0;
    #10.0; ADDR = 16'h81A9;
    #400.0; ADDR = 16'h81A8;
    #10.0; ADDR = 16'h81AA;
    #410.0; ADDR = 16'h81AB;
    #400.0; ADDR = 16'h81AC;
    #410.0; ADDR = 16'h1EC2;
    #490.0; ADDR = 16'h1EC3;
    #410.0; ADDR = 16'h81AD;
    #410.0; ADDR = 16'h81AE;
    #410.0; ADDR = 16'h81AF;
    #160.0; ADDR = 16'h1EA2;
    #10.0; ADDR = 16'h1EE2;
    #570.0; ADDR = 16'h1EE3;
    #400.0; ADDR = 16'h01AF;
    #10.0; ADDR = 16'h81AF;
    #400.0; ADDR = 16'h81A0;
    #10.0; ADDR = 16'h81B0;
    #650.0; ADDR = 16'h81A9;
    #410.0; ADDR = 16'h81AA;
    #410.0; ADDR = 16'h81AB;
    #400.0; ADDR = 16'h81A8;
    #10.0; ADDR = 16'h81AC;
    #400.0; ADDR = 16'h1880;
    #10.0; ADDR = 16'h1EC2;
    #490.0; ADDR = 16'h1EC3;
    #400.0; ADDR = 16'h00C3;
    #10.0; ADDR = 16'h81AD;
    #400.0; ADDR = 16'h81AC;
    #10.0; ADDR = 16'h81AE;
    #410.0; ADDR = 16'h81AF;
    #150.0; ADDR = 16'h80AF;
    #10.0; ADDR = 16'h1EE2;
    #570.0; ADDR = 16'h1EE3;
    #410.0; ADDR = 16'h81AF;
    #410.0; ADDR = 16'h81A0;
    #10.0; ADDR = 16'h81B0;
    #640.0; ADDR = 16'h81A0;
    #10.0; ADDR = 16'h81A9;
    #400.0; ADDR = 16'h81A8;
    #10.0; ADDR = 16'h81AA;
    #410.0; ADDR = 16'h81AB;
    #400.0; ADDR = 16'h81A8;
    #10.0; ADDR = 16'h81AC;
    #400.0; ADDR = 16'h1E80;
    #10.0; ADDR = 16'h1EC2;
    #490.0; ADDR = 16'h1EC3;
    #400.0; ADDR = 16'h01A9;
    #10.0; ADDR = 16'h81AD;
    #400.0; ADDR = 16'h81AC;
    #10.0; ADDR = 16'h81AE;
    #410.0; ADDR = 16'h81AF;
    #150.0; ADDR = 16'h98A3;
    #10.0; ADDR = 16'h1EE2;
    #570.0; ADDR = 16'h1EE3;
    #400.0; ADDR = 16'h06E3;
    #10.0; ADDR = 16'h81AF;
    #410.0; ADDR = 16'h81B0;
    #650.0; ADDR = 16'h81A0;
    #10.0; ADDR = 16'h81A9;
    #400.0; ADDR = 16'h81A8;
    #10.0; ADDR = 16'h81AA;
    #410.0; ADDR = 16'h81AB;
    #400.0; ADDR = 16'h81AC;
    #410.0; ADDR = 16'h1EC2;
    #490.0; ADDR = 16'h1EC3;
    #410.0; ADDR = 16'h81AD;
    #410.0; ADDR = 16'h81AC;
    #10.0; ADDR = 16'h81AE;
    #400.0; ADDR = 16'h81AF;
    #160.0; ADDR = 16'h1EA2;
    #10.0; ADDR = 16'h1EE2;
    #570.0; ADDR = 16'h1EE3;
    #400.0; ADDR = 16'h01AF;
    #10.0; ADDR = 16'h81AF;
    #400.0; ADDR = 16'h81A0;
    #10.0; ADDR = 16'h81B0;
    #650.0; ADDR = 16'h81A9;
    #410.0; ADDR = 16'h81AA;
    #410.0; ADDR = 16'h81AB;
    #400.0; ADDR = 16'h81A8;
    #10.0; ADDR = 16'h81AC;
    #400.0; ADDR = 16'h8880;
    #10.0; ADDR = 16'h1EC2;
    #490.0; ADDR = 16'h1EC3;
    #400.0; ADDR = 16'h00C3;
    #10.0; ADDR = 16'h81AD;
    #400.0; ADDR = 16'h81AC;
    #10.0; ADDR = 16'h81AE;
    #410.0; ADDR = 16'h81AF;
    #160.0; ADDR = 16'h1EE2;
    #570.0; ADDR = 16'h1EE3;
    #410.0; ADDR = 16'h81AF;
    #410.0; ADDR = 16'h81A0;
    #10.0; ADDR = 16'h81B0;
    #640.0; ADDR = 16'h81A0;
    #10.0; ADDR = 16'h81A9;
    #400.0; ADDR = 16'h81A8;
    #10.0; ADDR = 16'h81AA;
    #410.0; ADDR = 16'h81AB;
    #400.0; ADDR = 16'h81A8;
    #10.0; ADDR = 16'h81AC;
    #400.0; ADDR = 16'h1E80;
    #10.0; ADDR = 16'h1EC2;
    #490.0; ADDR = 16'h1EC3;
    #400.0; ADDR = 16'h01AD;
    #10.0; ADDR = 16'h81AD;
    #400.0; ADDR = 16'h81AC;
    #10.0; ADDR = 16'h81AE;
    #400.0; ADDR = 16'h1FAE;
    #10.0; ADDR = 16'h1FFF;
    #400.0; ADDR = 16'h1FFE;
    #410.0; ADDR = 16'h1FFD;
    #410.0; ADDR = 16'h1FFC;
    #410.0; ADDR = 16'h1FFB;
    #410.0; ADDR = 16'h1FFA;
    #410.0; ADDR = 16'h1FF9;
    #400.0; ADDR = 16'h1FF8;
    #410.0; ADDR = 16'h1FF0;
    #10.0; ADDR = 16'h1FF7;
    #400.0; ADDR = 16'h1FF6;
    #410.0; ADDR = 16'h1FF4;
    #10.0; ADDR = 16'h1FF5;
    #400.0; ADDR = 16'h1FF4;
    #410.0; ADDR = 16'hFFF0;
    #10.0; ADDR = 16'hFFF8;
    #410.0; ADDR = 16'hFFF9;
    #400.0; ADDR = 16'h81F5;
    #410.0; ADDR = 16'h81F6;
    #410.0; ADDR = 16'h81F7;
    #570.0; ADDR = 16'h082C;
    #490.0; ADDR = 16'h8168;
    #10.0; ADDR = 16'h81F8;
    #400.0; ADDR = 16'h81F9;
    #490.0; ADDR = 16'h81F8;
    #10.0; ADDR = 16'h81FA;
    #410.0; ADDR = 16'h81FB;
    #400.0; ADDR = 16'h81F8;
    #10.0; ADDR = 16'h81FC;
    #400.0; ADDR = 16'h81FD;
    #410.0; ADDR = 16'h7800;
    #820.0; ADDR = 16'h81FE;
    #410.0; ADDR = 16'h81FF;
    #490.0; ADDR = 16'h8200;
    #410.0; ADDR = 16'h8201;
    #410.0; ADDR = 16'h8202;
    #410.0; ADDR = 16'h8203;
    #400.0; ADDR = 16'h0200;
    #10.0; ADDR = 16'h5F84;
    #480.0; ADDR = 16'h0784;
    #10.0; ADDR = 16'h8204;
    #410.0; ADDR = 16'h8205;
    #490.0; ADDR = 16'h8206;
    #410.0; ADDR = 16'h8207;
    #240.0; ADDR = 16'h8208;
    #420.0; ADDR = 16'h8209;
    #400.0; ADDR = 16'h8208;
    #10.0; ADDR = 16'h820A;
    #410.0; ADDR = 16'h820B;
    #560.0; ADDR = 16'h0800;
    #10.0; ADDR = 16'h0834;
    #210.0; ADDR = 16'h0D34;
    #10.0; ADDR = 16'h0834;
    #340.0; ADDR = 16'h0034;
    #10.0; ADDR = 16'h820C;
    #410.0; ADDR = 16'h820D;
    #410.0; ADDR = 16'h820E;
    #570.0; ADDR = 16'h0808;
    #200.0; ADDR = 16'h0C08;
    #10.0; ADDR = 16'h0808;
    #280.0; ADDR = 16'h820F;
    #410.0; ADDR = 16'h8210;
    #250.0; ADDR = 16'h8211;
    #400.0; ADDR = 16'h8210;
    #10.0; ADDR = 16'h8212;
    #410.0; ADDR = 16'h8213;
    #560.0; ADDR = 16'h8813;
    #10.0; ADDR = 16'h0824;
    #480.0; ADDR = 16'h0024;
    #10.0; ADDR = 16'h8214;
    #410.0; ADDR = 16'h8215;
    #410.0; ADDR = 16'h8216;
    #570.0; ADDR = 16'h0824;
    #10.0; ADDR = 16'h0825;
    #560.0; ADDR = 16'h0005;
    #10.0; ADDR = 16'h8217;
    #400.0; ADDR = 16'h8218;
    #410.0; ADDR = 16'h8219;
    #570.0; ADDR = 16'h0801;
    #10.0; ADDR = 16'h0823;
    #480.0; ADDR = 16'h0023;
    #10.0; ADDR = 16'h821A;
    #400.0; ADDR = 16'h821B;
    #410.0; ADDR = 16'h821C;
    #570.0; ADDR = 16'h8814;
    #10.0; ADDR = 16'h0824;
    #570.0; ADDR = 16'h821D;
    #410.0; ADDR = 16'h821E;
    #420.0; ADDR = 16'h821F;
    #400.0; ADDR = 16'h8220;
    #400.0; ADDR = 16'h1200;
    #10.0; ADDR = 16'h5F81;
    #480.0; ADDR = 16'h0781;
    #10.0; ADDR = 16'h8221;
    #400.0; ADDR = 16'h8220;
    #10.0; ADDR = 16'h8222;
    #410.0; ADDR = 16'h8223;
    #490.0; ADDR = 16'h8224;
    #410.0; ADDR = 16'h8225;
    #400.0; ADDR = 16'h8224;
    #10.0; ADDR = 16'h8226;
    #410.0; ADDR = 16'h8227;
    #400.0; ADDR = 16'h8220;
    #10.0; ADDR = 16'h8228;
    #410.0; ADDR = 16'h8229;
    #400.0; ADDR = 16'h8228;
    #10.0; ADDR = 16'h822A;
    #410.0; ADDR = 16'h822B;
    #400.0; ADDR = 16'h8228;
    #10.0; ADDR = 16'h822C;
    #560.0; ADDR = 16'h0820;
    #10.0; ADDR = 16'h0823;
    #210.0; ADDR = 16'h0C23;
    #10.0; ADDR = 16'h0823;
    #340.0; ADDR = 16'h0023;
    #10.0; ADDR = 16'h822D;
    #410.0; ADDR = 16'h822E;
    #410.0; ADDR = 16'h822F;
    #400.0; ADDR = 16'h8221;
    #10.0; ADDR = 16'h8230;
    #400.0; ADDR = 16'h5A00;
    #10.0; ADDR = 16'h5F82;
    #480.0; ADDR = 16'h0782;
    #10.0; ADDR = 16'h8231;
    #400.0; ADDR = 16'h8230;
    #10.0; ADDR = 16'h8232;
    #410.0; ADDR = 16'h8233;
    #490.0; ADDR = 16'h8234;
    #410.0; ADDR = 16'h8235;
    #400.0; ADDR = 16'h8234;
    #10.0; ADDR = 16'h8236;
    #410.0; ADDR = 16'h8237;
    #400.0; ADDR = 16'h8230;
    #10.0; ADDR = 16'h8238;
    #410.0; ADDR = 16'h8239;
    #400.0; ADDR = 16'h8238;
    #10.0; ADDR = 16'h823A;
    #410.0; ADDR = 16'h823B;
    #560.0; ADDR = 16'h0823;
    #570.0; ADDR = 16'h0023;
    #10.0; ADDR = 16'h823C;
    #410.0; ADDR = 16'h823D;
    #400.0; ADDR = 16'h823C;
    #10.0; ADDR = 16'h823E;
    #570.0; ADDR = 16'h0823;
    #570.0; ADDR = 16'h823F;
    #410.0; ADDR = 16'h8240;
    #410.0; ADDR = 16'h8241;
    #410.0; ADDR = 16'h8242;
    #400.0; ADDR = 16'h8200;
    #10.0; ADDR = 16'h5F80;
    #490.0; ADDR = 16'h8243;
    #410.0; ADDR = 16'h8244;
    #410.0; ADDR = 16'h8245;
    #490.0; ADDR = 16'h8246;
    #410.0; ADDR = 16'h8247;
    #400.0; ADDR = 16'h8241;
    #10.0; ADDR = 16'h8248;
    #570.0; ADDR = 16'h0823;
    #570.0; ADDR = 16'h0001;
    #10.0; ADDR = 16'h8249;
    #400.0; ADDR = 16'h824B;
    #10.0; ADDR = 16'h824A;
    #400.0; ADDR = 16'h824B;
    #570.0; ADDR = 16'h0803;
    #10.0; ADDR = 16'h0823;
    #210.0; ADDR = 16'h0C23;
    #10.0; ADDR = 16'h0823;
    #340.0; ADDR = 16'h0023;
    #10.0; ADDR = 16'h824C;
    #410.0; ADDR = 16'h824D;
    #410.0; ADDR = 16'h824E;
    #570.0; ADDR = 16'h081A;
    #200.0; ADDR = 16'h0C1A;
    #10.0; ADDR = 16'h081A;
    #280.0; ADDR = 16'h824F;
    #410.0; ADDR = 16'h9250;
    #10.0; ADDR = 16'h8250;
    #650.0; ADDR = 16'h8269;
    #400.0; ADDR = 16'h8268;
    #10.0; ADDR = 16'h826A;
    #410.0; ADDR = 16'h826B;
    #560.0; ADDR = 16'h806B;
    #10.0; ADDR = 16'h0819;
    #200.0; ADDR = 16'h1B19;
    #10.0; ADDR = 16'h0819;
    #270.0; ADDR = 16'h0019;
    #10.0; ADDR = 16'h826C;
    #410.0; ADDR = 16'h826D;
    #650.0; ADDR = 16'h8200;
    #10.0; ADDR = 16'h8282;
    #410.0; ADDR = 16'h8283;
    #400.0; ADDR = 16'h8284;
    #570.0; ADDR = 16'h0804;
    #10.0; ADDR = 16'h081F;
    #480.0; ADDR = 16'h0007;
    #10.0; ADDR = 16'h8285;
    #400.0; ADDR = 16'h8287;
    #10.0; ADDR = 16'h8286;
    #650.0; ADDR = 16'h829F;
    #410.0; ADDR = 16'h82A0;
    #410.0; ADDR = 16'h82A1;
    #570.0; ADDR = 16'h081E;
    #490.0; ADDR = 16'h82A2;
    #410.0; ADDR = 16'h82A3;
    #650.0; ADDR = 16'h82A1;
    #10.0; ADDR = 16'h82B8;
    #410.0; ADDR = 16'h82B9;
    #400.0; ADDR = 16'h82B8;
    #10.0; ADDR = 16'h82BA;
    #560.0; ADDR = 16'h88BA;
    #10.0; ADDR = 16'h0823;
    #480.0; ADDR = 16'h0023;
    #10.0; ADDR = 16'h82BB;
    #410.0; ADDR = 16'h82BC;
    #410.0; ADDR = 16'h82BD;
    #570.0; ADDR = 16'h0824;
    #570.0; ADDR = 16'h0024;
    #10.0; ADDR = 16'h82BE;
    #400.0; ADDR = 16'h82BF;
    #410.0; ADDR = 16'h82C0;
    #420.0; ADDR = 16'h82C1;
    #560.0; ADDR = 16'h0801;
    #10.0; ADDR = 16'h0825;
    #560.0; ADDR = 16'h0025;
    #10.0; ADDR = 16'h82C2;
    #410.0; ADDR = 16'h82C3;
    #490.0; ADDR = 16'h82C4;
    #410.0; ADDR = 16'h82C5;
    #650.0; ADDR = 16'h8340;
    #410.0; ADDR = 16'h8341;
    #410.0; ADDR = 16'h8342;
    #570.0; ADDR = 16'h0814;
    #10.0; ADDR = 16'h0834;
    #480.0; ADDR = 16'h0100;
    #10.0; ADDR = 16'h8343;
    #400.0; ADDR = 16'h8347;
    #10.0; ADDR = 16'h8344;
    #650.0; ADDR = 16'h834A;
    #410.0; ADDR = 16'h834B;
    #410.0; ADDR = 16'h834C;
    #410.0; ADDR = 16'h834D;
    #400.0; ADDR = 16'h1A00;
    #10.0; ADDR = 16'h1E82;
    #490.0; ADDR = 16'h1E83;
    #400.0; ADDR = 16'h0783;
    #10.0; ADDR = 16'h834E;
    #410.0; ADDR = 16'h834F;
    #400.0; ADDR = 16'h8350;
    #420.0; ADDR = 16'h8351;
    #400.0; ADDR = 16'h1E00;
    #10.0; ADDR = 16'h1E80;
    #490.0; ADDR = 16'h1E81;
    #400.0; ADDR = 16'h0352;
    #10.0; ADDR = 16'h8352;
    #400.0; ADDR = 16'h8353;
    #660.0; ADDR = 16'h8366;
    #410.0; ADDR = 16'h8367;
    #400.0; ADDR = 16'h8360;
    #10.0; ADDR = 16'h8368;
    #570.0; ADDR = 16'h0801;
    #480.0; ADDR = 16'h0001;
    #10.0; ADDR = 16'h8369;
    #410.0; ADDR = 16'h836A;
    #650.0; ADDR = 16'h8302;
    #10.0; ADDR = 16'h8385;
    #400.0; ADDR = 16'h8384;
    #10.0; ADDR = 16'h8386;
    #410.0; ADDR = 16'h8387;
    #400.0; ADDR = 16'h8388;
    #410.0; ADDR = 16'h5F88;
    #490.0; ADDR = 16'h0389;
    #10.0; ADDR = 16'h8389;
    #400.0; ADDR = 16'h8388;
    #10.0; ADDR = 16'h838A;
    #400.0; ADDR = 16'h838B;
    #570.0; ADDR = 16'h0806;
    #900.0; ADDR = 16'h0004;
    #10.0; ADDR = 16'h838C;
    #410.0; ADDR = 16'h838D;
    #480.0; ADDR = 16'h838C;
    #10.0; ADDR = 16'h838E;
    #410.0; ADDR = 16'h838F;
    #400.0; ADDR = 16'h8380;
    #10.0; ADDR = 16'h8390;
    #560.0; ADDR = 16'h8890;
    #10.0; ADDR = 16'h0801;
    #570.0; ADDR = 16'h8391;
    #410.0; ADDR = 16'h8392;
    #410.0; ADDR = 16'h8393;
    #570.0; ADDR = 16'h083A;
    #500.0; ADDR = 16'h083B;
    #400.0; ADDR = 16'h8310;
    #10.0; ADDR = 16'h8394;
    #410.0; ADDR = 16'h8395;
    #400.0; ADDR = 16'h8394;
    #10.0; ADDR = 16'h8396;
    #490.0; ADDR = 16'h8397;
    #400.0; ADDR = 16'h8390;
    #10.0; ADDR = 16'h8398;
    #490.0; ADDR = 16'h8399;
    #400.0; ADDR = 16'h8398;
    #10.0; ADDR = 16'h839A;
    #410.0; ADDR = 16'h839B;
    #400.0; ADDR = 16'h839C;
    #420.0; ADDR = 16'h839D;
    #400.0; ADDR = 16'h839E;
    #400.0; ADDR = 16'h829E;
    #10.0; ADDR = 16'h5A00;
    #660.0; ADDR = 16'h5A01;
    #640.0; ADDR = 16'h0201;
    #10.0; ADDR = 16'h839F;
    #410.0; ADDR = 16'h83A0;
    #410.0; ADDR = 16'h83A1;
    #570.0; ADDR = 16'h083C;
    #490.0; ADDR = 16'h083D;
    #120.0; ADDR = 16'h0C3D;
    #10.0; ADDR = 16'h083D;
    #280.0; ADDR = 16'h83A0;
    #10.0; ADDR = 16'h83A2;
    #410.0; ADDR = 16'h83A3;
    #400.0; ADDR = 16'h83A0;
    #10.0; ADDR = 16'h83A4;
    #490.0; ADDR = 16'h83A5;
    #400.0; ADDR = 16'h83A4;
    #10.0; ADDR = 16'h83A6;
    #490.0; ADDR = 16'h83A7;
    #400.0; ADDR = 16'h83A8;
    #410.0; ADDR = 16'h83A9;
    #410.0; ADDR = 16'h83AA;
    #420.0; ADDR = 16'h83AB;
    #400.0; ADDR = 16'h83AC;
    #400.0; ADDR = 16'h82AC;
    #10.0; ADDR = 16'h7A00;
    #900.0; ADDR = 16'h7A01;
    #650.0; ADDR = 16'h0201;
    #10.0; ADDR = 16'h83AD;
    #400.0; ADDR = 16'h83AE;
    #410.0; ADDR = 16'h83AF;
    #570.0; ADDR = 16'h88AF;
    #10.0; ADDR = 16'h083E;
    #490.0; ADDR = 16'h083F;
    #400.0; ADDR = 16'h0031;
    #10.0; ADDR = 16'h83B0;
    #400.0; ADDR = 16'h83B1;
    #410.0; ADDR = 16'h83B3;
    #10.0; ADDR = 16'h83B2;
    #410.0; ADDR = 16'h83B3;
    #400.0; ADDR = 16'h5800;
    #10.0; ADDR = 16'h580C;
    #640.0; ADDR = 16'h000C;
    #10.0; ADDR = 16'h83B4;
    #410.0; ADDR = 16'h83B5;
    #410.0; ADDR = 16'h83B6;
    #410.0; ADDR = 16'h83B7;
    #400.0; ADDR = 16'h6004;
    #10.0; ADDR = 16'h780C;
    #650.0; ADDR = 16'h03B8;
    #10.0; ADDR = 16'h83B8;
    #400.0; ADDR = 16'h83B9;
    #410.0; ADDR = 16'h83BA;
    #570.0; ADDR = 16'h0808;
    #490.0; ADDR = 16'h0008;
    #10.0; ADDR = 16'h83BB;
    #400.0; ADDR = 16'h83BF;
    #10.0; ADDR = 16'h83BC;
    #410.0; ADDR = 16'h83BD;
    #400.0; ADDR = 16'h83BC;
    #10.0; ADDR = 16'h83BE;
    #240.0; ADDR = 16'h83BF;
    #410.0; ADDR = 16'h83C0;
    #410.0; ADDR = 16'h83C1;
    #570.0; ADDR = 16'h0809;
    #490.0; ADDR = 16'h83C0;
    #10.0; ADDR = 16'h83C2;
    #400.0; ADDR = 16'h83C3;
    #410.0; ADDR = 16'h83C4;
    #410.0; ADDR = 16'h83C5;
    #240.0; ADDR = 16'h83C4;
    #10.0; ADDR = 16'h83C6;
    #410.0; ADDR = 16'h83C7;
    #400.0; ADDR = 16'h83C0;
    #10.0; ADDR = 16'h83C8;
    #560.0; ADDR = 16'h88C8;
    #10.0; ADDR = 16'h080A;
    #200.0; ADDR = 16'h0C0A;
    #10.0; ADDR = 16'h080A;
    #270.0; ADDR = 16'h000A;
    #10.0; ADDR = 16'h83C9;
    #410.0; ADDR = 16'h83CA;
    #410.0; ADDR = 16'h83CB;
    #400.0; ADDR = 16'h83C8;
    #10.0; ADDR = 16'h83CC;
    #250.0; ADDR = 16'h83CD;
    #400.0; ADDR = 16'h83CE;
    #490.0; ADDR = 16'h83CF;
    #410.0; ADDR = 16'h83C0;
    #10.0; ADDR = 16'h83D0;
    #410.0; ADDR = 16'h83D1;
    #400.0; ADDR = 16'h83D2;
    #410.0; ADDR = 16'h0927;
    #900.0; ADDR = 16'h83D3;
    #410.0; ADDR = 16'h83D4;
    #650.0; ADDR = 16'h83D0;
    #10.0; ADDR = 16'h83D8;
    #410.0; ADDR = 16'h83D9;
    #400.0; ADDR = 16'h83D8;
    #10.0; ADDR = 16'h83DA;
    #560.0; ADDR = 16'h88DA;
    #10.0; ADDR = 16'h0826;
    #190.0; ADDR = 16'h0C26;
    #10.0; ADDR = 16'h0826;
    #290.0; ADDR = 16'h0827;
    #400.0; ADDR = 16'h0003;
    #10.0; ADDR = 16'h83DB;
    #410.0; ADDR = 16'h83DC;
    #410.0; ADDR = 16'h83DD;
    #560.0; ADDR = 16'h8BDD;
    #10.0; ADDR = 16'h0827;
    #570.0; ADDR = 16'h0828;
    #410.0; ADDR = 16'h83DE;
    #410.0; ADDR = 16'h83DF;
    #410.0; ADDR = 16'h83E0;
    #410.0; ADDR = 16'h83E1;
    #400.0; ADDR = 16'h81E1;
    #10.0; ADDR = 16'h0926;
    #480.0; ADDR = 16'h0126;
    #10.0; ADDR = 16'h83E2;
    #410.0; ADDR = 16'h83E3;
    #410.0; ADDR = 16'h83E4;
    #570.0; ADDR = 16'h0826;
    #570.0; ADDR = 16'h0024;
    #10.0; ADDR = 16'h83E5;
    #400.0; ADDR = 16'h83E7;
    #10.0; ADDR = 16'h83E6;
    #410.0; ADDR = 16'h83E7;
    #400.0; ADDR = 16'h83E0;
    #10.0; ADDR = 16'h83E8;
    #400.0; ADDR = 16'h0929;
    #900.0; ADDR = 16'h83E9;
    #410.0; ADDR = 16'h83EA;
    #660.0; ADDR = 16'h83EE;
    #410.0; ADDR = 16'h83EF;
    #400.0; ADDR = 16'h83E0;
    #10.0; ADDR = 16'h83F0;
    #560.0; ADDR = 16'h8AF0;
    #10.0; ADDR = 16'h0829;
    #490.0; ADDR = 16'h082A;
    #120.0; ADDR = 16'h382A;
    #10.0; ADDR = 16'h082A;
    #270.0; ADDR = 16'h0022;
    #10.0; ADDR = 16'h83F1;
    #410.0; ADDR = 16'h83F2;
    #410.0; ADDR = 16'h83F3;
    #570.0; ADDR = 16'h082A;
    #570.0; ADDR = 16'h082B;
    #410.0; ADDR = 16'h83F4;
    #410.0; ADDR = 16'h83F5;
    #410.0; ADDR = 16'h83F4;
    #10.0; ADDR = 16'h83F6;
    #400.0; ADDR = 16'h83F7;
    #410.0; ADDR = 16'h0928;
    #200.0; ADDR = 16'h1D28;
    #10.0; ADDR = 16'h0928;
    #270.0; ADDR = 16'h0128;
    #10.0; ADDR = 16'h83F8;
    #410.0; ADDR = 16'h83F9;
    #410.0; ADDR = 16'h83FA;
    #570.0; ADDR = 16'h0829;
    #220.0; ADDR = 16'h1829;
    #10.0; ADDR = 16'h0829;
    #340.0; ADDR = 16'h0029;
    #10.0; ADDR = 16'h83FB;
    #400.0; ADDR = 16'h83FE;
    #10.0; ADDR = 16'h83FC;
    #650.0; ADDR = 16'h8419;
    #410.0; ADDR = 16'h841A;
    #410.0; ADDR = 16'h841B;
    #570.0; ADDR = 16'h082C;
    #490.0; ADDR = 16'h841C;
    #410.0; ADDR = 16'h841D;
    #410.0; ADDR = 16'h841E;
    #410.0; ADDR = 16'h841F;
    #400.0; ADDR = 16'h8017;
    #10.0; ADDR = 16'h7800;
    #650.0; ADDR = 16'h0420;
    #10.0; ADDR = 16'h8420;
    #400.0; ADDR = 16'h8421;
    #410.0; ADDR = 16'h8422;
    #570.0; ADDR = 16'h0800;
    #10.0; ADDR = 16'h0808;
    #480.0; ADDR = 16'h0000;
    #10.0; ADDR = 16'h8423;
    #400.0; ADDR = 16'h8427;
    #10.0; ADDR = 16'h8424;
    #400.0; ADDR = 16'h8425;
    #410.0; ADDR = 16'h8424;
    #10.0; ADDR = 16'h8426;
    #410.0; ADDR = 16'h8427;
    #400.0; ADDR = 16'h8420;
    #10.0; ADDR = 16'h8428;
    #400.0; ADDR = 16'h8429;
    #160.0; ADDR = 16'hE409;
    #10.0; ADDR = 16'hE44F;
    #240.0; ADDR = 16'hE451;
    #410.0; ADDR = 16'hE452;
    #400.0; ADDR = 16'h8052;
    #10.0; ADDR = 16'h8AA7;
    #160.0; ADDR = 16'h1BA3;
    #10.0; ADDR = 16'h1FF3;
    #400.0; ADDR = 16'h1FF2;
    #410.0; ADDR = 16'h8AA7;
    #410.0; ADDR = 16'h8AA8;
    #410.0; ADDR = 16'h8AA9;
    #570.0; ADDR = 16'h0802;
    #500.0; ADDR = 16'h8AAA;
    #400.0; ADDR = 16'h8AAB;
    #410.0; ADDR = 16'h8AAC;
    #490.0; ADDR = 16'h8B84;
    #10.0; ADDR = 16'h8B85;
    #400.0; ADDR = 16'h8B84;
    #10.0; ADDR = 16'h8B86;
    #410.0; ADDR = 16'h8B87;
    #560.0; ADDR = 16'h0809;
    #500.0; ADDR = 16'h8B88;
    #400.0; ADDR = 16'h8B89;
    #410.0; ADDR = 16'h8B88;
    #10.0; ADDR = 16'h8B8A;
    #400.0; ADDR = 16'h8B8B;
    #410.0; ADDR = 16'h8B88;
    #10.0; ADDR = 16'h8B8C;
    #410.0; ADDR = 16'h8B8D;
    #400.0; ADDR = 16'h8B8C;
    #10.0; ADDR = 16'h8B8E;
    #150.0; ADDR = 16'hE08E;
    #10.0; ADDR = 16'hE4E0;
    #240.0; ADDR = 16'hE4E6;
    #420.0; ADDR = 16'hE4E7;
    #400.0; ADDR = 16'h8DD5;
    #410.0; ADDR = 16'h8DD6;
    #410.0; ADDR = 16'h8DD7;
    #570.0; ADDR = 16'h080A;
    #490.0; ADDR = 16'h0908;
    #10.0; ADDR = 16'h8DD8;
    #400.0; ADDR = 16'h8DD9;
    #410.0; ADDR = 16'h8DDA;
    #410.0; ADDR = 16'h8DDB;
    #410.0; ADDR = 16'h8DD8;
    #10.0; ADDR = 16'h8DDC;
    #400.0; ADDR = 16'h8DDD;
    #410.0; ADDR = 16'h8DDE;
    #160.0; ADDR = 16'hE502;
    #250.0; ADDR = 16'hE506;
    #410.0; ADDR = 16'hE507;
    #400.0; ADDR = 16'h8407;
    #10.0; ADDR = 16'h8E69;
    #400.0; ADDR = 16'h8E68;
    #10.0; ADDR = 16'h8E6A;
    #410.0; ADDR = 16'h8E6B;
    #570.0; ADDR = 16'h0829;
    #490.0; ADDR = 16'h8E6C;
    #410.0; ADDR = 16'h8E6D;
    #490.0; ADDR = 16'h8E6C;
    #10.0; ADDR = 16'h8E6E;
    #400.0; ADDR = 16'h8E6F;
    #650.0; ADDR = 16'h8E2B;
    #10.0; ADDR = 16'h8EAA;
    #410.0; ADDR = 16'h8EAB;
    #400.0; ADDR = 16'h8EA8;
    #10.0; ADDR = 16'h8EAC;
    #560.0; ADDR = 16'h88AC;
    #10.0; ADDR = 16'h0806;
    #490.0; ADDR = 16'h8EAD;
    #410.0; ADDR = 16'h8EAE;
    #490.0; ADDR = 16'h8EAF;
    #410.0; ADDR = 16'h8EB0;
    #250.0; ADDR = 16'h8EB1;
    #400.0; ADDR = 16'h8EB0;
    #10.0; ADDR = 16'h8EB2;
    #490.0; ADDR = 16'h8EB3;
    #400.0; ADDR = 16'h8EB0;
    #10.0; ADDR = 16'h8EB4;
    #640.0; ADDR = 16'h9EB4;
    #10.0; ADDR = 16'h1FF1;
    #410.0; ADDR = 16'h1FF0;
    #400.0; ADDR = 16'h0FF0;
    #10.0; ADDR = 16'h8F14;
    #410.0; ADDR = 16'h8F15;
    #400.0; ADDR = 16'h8F14;
    #10.0; ADDR = 16'h8F16;
    #410.0; ADDR = 16'h8F17;
    #400.0; ADDR = 16'h8F10;
    #10.0; ADDR = 16'h8F18;
    #410.0; ADDR = 16'h8F19;
    #400.0; ADDR = 16'h8F18;
    #10.0; ADDR = 16'h8F1A;
    #400.0; ADDR = 16'h8F1B;
    #410.0; ADDR = 16'h8F1C;
    #160.0; ADDR = 16'hE508;
    #570.0; ADDR = 16'h8D08;
    #10.0; ADDR = 16'h8F1C;
    #410.0; ADDR = 16'h8F1D;
    #240.0; ADDR = 16'h8F1C;
    #10.0; ADDR = 16'h8F1E;
    #400.0; ADDR = 16'h8F1F;
    #410.0; ADDR = 16'h8F20;
    #410.0; ADDR = 16'h8F21;
    #240.0; ADDR = 16'h8F20;
    #10.0; ADDR = 16'h8F22;
    #410.0; ADDR = 16'h8F23;
    #400.0; ADDR = 16'h8F20;
    #10.0; ADDR = 16'h8F24;
    #410.0; ADDR = 16'h8F25;
    #480.0; ADDR = 16'h6419;
    #820.0; ADDR = 16'h8F06;
    #10.0; ADDR = 16'h8F26;
    #400.0; ADDR = 16'h8F27;
    #410.0; ADDR = 16'h8F28;
    #160.0; ADDR = 16'hE508;
    #10.0; ADDR = 16'hE509;
    #560.0; ADDR = 16'h8D09;
    #10.0; ADDR = 16'h8F28;
    #410.0; ADDR = 16'h8F29;
    #400.0; ADDR = 16'h8F28;
    #10.0; ADDR = 16'h8F2A;
    #410.0; ADDR = 16'h8F2B;
    #480.0; ADDR = 16'hE42B;
    #10.0; ADDR = 16'h6459;
    #650.0; ADDR = 16'h8F2C;
    #410.0; ADDR = 16'h8F2D;
    #410.0; ADDR = 16'h8F2E;
    #730.0; ADDR = 16'h442A;
    #10.0; ADDR = 16'h4459;
    #730.0; ADDR = 16'h8F0F;
    #10.0; ADDR = 16'h8F2F;
    #400.0; ADDR = 16'h8F30;
    #410.0; ADDR = 16'h8F31;
    #160.0; ADDR = 16'h4419;
    #980.0; ADDR = 16'h0C11;
    #10.0; ADDR = 16'h8F31;
    #400.0; ADDR = 16'h8F33;
    #10.0; ADDR = 16'h8F32;
    #650.0; ADDR = 16'h8F1A;
    #410.0; ADDR = 16'h8F1B;
    #400.0; ADDR = 16'h8F19;
    #10.0; ADDR = 16'h8F1C;
    #160.0; ADDR = 16'hE508;
    #10.0; ADDR = 16'hE50A;
    #560.0; ADDR = 16'h8D08;
    #10.0; ADDR = 16'h8F1C;
    #410.0; ADDR = 16'h8F1D;
    #650.0; ADDR = 16'h8F33;
    #410.0; ADDR = 16'h8F34;
    #410.0; ADDR = 16'h8F35;
    #730.0; ADDR = 16'h441B;
    #330.0; ADDR = 16'h8F32;
    #10.0; ADDR = 16'h8F36;
    #400.0; ADDR = 16'h8F37;
    #650.0; ADDR = 16'h8F12;
    #10.0; ADDR = 16'h8F1A;
    #410.0; ADDR = 16'h8F1B;
    #400.0; ADDR = 16'h8F18;
    #10.0; ADDR = 16'h8F1C;
    #150.0; ADDR = 16'hE50C;
    #10.0; ADDR = 16'hE50B;
    #570.0; ADDR = 16'h8F1C;
    #410.0; ADDR = 16'h8F1D;
    #240.0; ADDR = 16'h8F1C;
    #10.0; ADDR = 16'h8F1E;
    #410.0; ADDR = 16'h8F1F;
    #400.0; ADDR = 16'h8F20;
    #420.0; ADDR = 16'h8F21;
    #240.0; ADDR = 16'h8F22;
    #410.0; ADDR = 16'h8F23;
    #400.0; ADDR = 16'h8F20;
    #10.0; ADDR = 16'h8F24;
    #410.0; ADDR = 16'h8F25;
    #480.0; ADDR = 16'hE525;
    #10.0; ADDR = 16'h641B;
    #730.0; ADDR = 16'h0F02;
    #10.0; ADDR = 16'h8F26;
    #400.0; ADDR = 16'h8F27;
    #410.0; ADDR = 16'h8F28;
    #160.0; ADDR = 16'hE508;
    #10.0; ADDR = 16'hE50C;
    #560.0; ADDR = 16'hC50C;
    #10.0; ADDR = 16'h8F28;
    #410.0; ADDR = 16'h8F29;
    #400.0; ADDR = 16'h8F28;
    #10.0; ADDR = 16'h8F2A;
    #410.0; ADDR = 16'h8F2B;
    #480.0; ADDR = 16'hE42B;
    #10.0; ADDR = 16'h645B;
    #650.0; ADDR = 16'h8F0C;
    #10.0; ADDR = 16'h8F2C;
    #400.0; ADDR = 16'h8F2D;
    #410.0; ADDR = 16'h8F2E;
    #730.0; ADDR = 16'hC42A;
    #10.0; ADDR = 16'h445B;
    #730.0; ADDR = 16'h8F0B;
    #10.0; ADDR = 16'h8F2F;
    #400.0; ADDR = 16'h8F30;
    #410.0; ADDR = 16'h8F31;
    #160.0; ADDR = 16'h4411;
    #10.0; ADDR = 16'h441B;
    #970.0; ADDR = 16'h0C11;
    #10.0; ADDR = 16'h8F31;
    #410.0; ADDR = 16'h8F32;
    #650.0; ADDR = 16'h8F1A;
    #410.0; ADDR = 16'h8F1B;
    #410.0; ADDR = 16'h8F1C;
    #160.0; ADDR = 16'hE50C;
    #10.0; ADDR = 16'hE50D;
    #560.0; ADDR = 16'h8D0C;
    #10.0; ADDR = 16'h8F1C;
    #410.0; ADDR = 16'h8F1D;
    #650.0; ADDR = 16'h8F33;
    #410.0; ADDR = 16'h8F34;
    #410.0; ADDR = 16'h8F35;
    #730.0; ADDR = 16'h441D;
    #330.0; ADDR = 16'h8F16;
    #10.0; ADDR = 16'h8F36;
    #400.0; ADDR = 16'h8F37;
    #650.0; ADDR = 16'h8F12;
    #10.0; ADDR = 16'h8F1A;
    #410.0; ADDR = 16'h8F1B;
    #400.0; ADDR = 16'h8F18;
    #10.0; ADDR = 16'h8F1C;
    #150.0; ADDR = 16'hE50C;
    #10.0; ADDR = 16'hE50E;
    #560.0; ADDR = 16'h850E;
    #10.0; ADDR = 16'h8F1C;
    #410.0; ADDR = 16'h8F1D;
    #240.0; ADDR = 16'h8F1C;
    #10.0; ADDR = 16'h8F1E;
    #410.0; ADDR = 16'h8F1F;
    #400.0; ADDR = 16'h8F20;
    #410.0; ADDR = 16'h8F21;
    #250.0; ADDR = 16'h8F22;
    #410.0; ADDR = 16'h8F23;
    #400.0; ADDR = 16'h8F20;
    #10.0; ADDR = 16'h8F24;
    #410.0; ADDR = 16'h8F25;
    #480.0; ADDR = 16'h640D;
    #10.0; ADDR = 16'h641D;
    #730.0; ADDR = 16'h8F06;
    #10.0; ADDR = 16'h8F26;
    #400.0; ADDR = 16'h8F27;
    #410.0; ADDR = 16'h8F28;
    #160.0; ADDR = 16'hE50E;
    #10.0; ADDR = 16'hE50F;
    #560.0; ADDR = 16'h8D0B;
    #10.0; ADDR = 16'h8F28;
    #410.0; ADDR = 16'h8F29;
    #400.0; ADDR = 16'h8F28;
    #10.0; ADDR = 16'h8F2A;
    #410.0; ADDR = 16'h8F2B;
    #480.0; ADDR = 16'hE42B;
    #10.0; ADDR = 16'h645D;
    #650.0; ADDR = 16'h8F0C;
    #10.0; ADDR = 16'h8F2C;
    #400.0; ADDR = 16'h8F2D;
    #410.0; ADDR = 16'h8F2E;
    #730.0; ADDR = 16'hC42E;
    #10.0; ADDR = 16'h445D;
    #730.0; ADDR = 16'h8F0D;
    #10.0; ADDR = 16'h8F2F;
    #400.0; ADDR = 16'h8F30;
    #410.0; ADDR = 16'h8F31;
    #160.0; ADDR = 16'h4415;
    #10.0; ADDR = 16'h441D;
    #970.0; ADDR = 16'h0C11;
    #10.0; ADDR = 16'h8F31;
    #410.0; ADDR = 16'h8F32;
    #650.0; ADDR = 16'h8F1A;
    #410.0; ADDR = 16'h8F1B;
    #410.0; ADDR = 16'h8F1C;
    #160.0; ADDR = 16'hE510;
    #570.0; ADDR = 16'h8510;
    #10.0; ADDR = 16'h8F1C;
    #410.0; ADDR = 16'h8F1D;
    #650.0; ADDR = 16'h8F33;
    #410.0; ADDR = 16'h8F34;
    #410.0; ADDR = 16'h8F35;
    #730.0; ADDR = 16'h441F;
    #330.0; ADDR = 16'h8F16;
    #10.0; ADDR = 16'h8F36;
    #400.0; ADDR = 16'h8F37;
    #650.0; ADDR = 16'h8F12;
    #10.0; ADDR = 16'h8F1A;
    #410.0; ADDR = 16'h8F1B;
    #400.0; ADDR = 16'h8F18;
    #10.0; ADDR = 16'h8F1C;
    #150.0; ADDR = 16'hE514;
    #10.0; ADDR = 16'hE511;
    #560.0; ADDR = 16'hC511;
    #10.0; ADDR = 16'h8F1C;
    #410.0; ADDR = 16'h8F1D;
    #240.0; ADDR = 16'h8F1C;
    #10.0; ADDR = 16'h8F1E;
    #410.0; ADDR = 16'h8F1F;
    #400.0; ADDR = 16'h8F20;
    #410.0; ADDR = 16'h8F21;
    #250.0; ADDR = 16'h8F22;
    #410.0; ADDR = 16'h8F23;
    #400.0; ADDR = 16'h8F20;
    #10.0; ADDR = 16'h8F24;
    #410.0; ADDR = 16'h8F25;
    #480.0; ADDR = 16'h640D;
    #10.0; ADDR = 16'h641F;
    #730.0; ADDR = 16'h8F06;
    #10.0; ADDR = 16'h8F26;
    #400.0; ADDR = 16'h8F27;
    #410.0; ADDR = 16'h8F28;
    #160.0; ADDR = 16'hE500;
    #10.0; ADDR = 16'hE512;
    #560.0; ADDR = 16'h8D00;
    #10.0; ADDR = 16'h8F28;
    #410.0; ADDR = 16'h8F29;
    #400.0; ADDR = 16'h8F28;
    #10.0; ADDR = 16'h8F2A;
    #410.0; ADDR = 16'h8F2B;
    #480.0; ADDR = 16'hE40B;
    #10.0; ADDR = 16'h645F;
    #650.0; ADDR = 16'h8F2C;
    #410.0; ADDR = 16'h8F2D;
    #410.0; ADDR = 16'h8F2E;
    #730.0; ADDR = 16'h440E;
    #10.0; ADDR = 16'h445F;
    #730.0; ADDR = 16'h8F0F;
    #10.0; ADDR = 16'h8F2F;
    #400.0; ADDR = 16'h8F30;
    #410.0; ADDR = 16'h8F31;
    #160.0; ADDR = 16'h4417;
    #10.0; ADDR = 16'h441F;

end
initial
begin
    DATA = 8'hFF;
    #560.0; DATA = 8'h75;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'hF8;
    #330.0; DATA = 8'hFF;
    #330.0; DATA = 8'h43;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h07;
    #320.0; DATA = 8'h0F;
    #10.0; DATA = 8'hFF;
    #80.0; DATA = 8'h1E;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'hC2;
    #320.0; DATA = 8'hFF;
    #200.0; DATA = 8'h9E;
    #10.0; DATA = 8'h1E;
    #380.0; DATA = 8'hDE;
    #20.0; DATA = 8'hFA;
    #10.0; DATA = 8'hE2;
    #370.0; DATA = 8'h41;
    #320.0; DATA = 8'hE2;
    #80.0; DATA = 8'hA2;
    #10.0; DATA = 8'h26;
    #320.0; DATA = 8'hE2;
    #10.0; DATA = 8'hEB;
    #10.0; DATA = 8'hEF;
    #400.0; DATA = 8'hFF;
    #20.0; DATA = 8'hFA;
    #10.0; DATA = 8'hFF;
    #780.0; DATA = 8'h75;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hF8;
    #330.0; DATA = 8'hFF;
    #320.0; DATA = 8'hF7;
    #10.0; DATA = 8'h43;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'h07;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h1E;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hC2;
    #330.0; DATA = 8'hFF;
    #190.0; DATA = 8'hFE;
    #10.0; DATA = 8'h1E;
    #390.0; DATA = 8'hDE;
    #20.0; DATA = 8'hF2;
    #10.0; DATA = 8'hE2;
    #360.0; DATA = 8'h41;
    #330.0; DATA = 8'hE2;
    #80.0; DATA = 8'h26;
    #330.0; DATA = 8'hE2;
    #10.0; DATA = 8'hEF;
    #410.0; DATA = 8'hFF;
    #10.0; DATA = 8'hFA;
    #10.0; DATA = 8'hFE;
    #10.0; DATA = 8'hFF;
    #780.0; DATA = 8'h75;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'hF8;
    #320.0; DATA = 8'hFF;
    #330.0; DATA = 8'h43;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h07;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h1E;
    #320.0; DATA = 8'h1F;
    #10.0; DATA = 8'hFF;
    #80.0; DATA = 8'hC2;
    #320.0; DATA = 8'hC3;
    #10.0; DATA = 8'hFF;
    #190.0; DATA = 8'hDE;
    #10.0; DATA = 8'h1E;
    #380.0; DATA = 8'hDE;
    #20.0; DATA = 8'hFA;
    #10.0; DATA = 8'hE2;
    #370.0; DATA = 8'h41;
    #320.0; DATA = 8'h42;
    #10.0; DATA = 8'hE2;
    #80.0; DATA = 8'h26;
    #320.0; DATA = 8'hE2;
    #10.0; DATA = 8'hE3;
    #10.0; DATA = 8'hEB;
    #400.0; DATA = 8'hFF;
    #20.0; DATA = 8'hFA;
    #10.0; DATA = 8'hFF;
    #780.0; DATA = 8'h75;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hF8;
    #330.0; DATA = 8'hFF;
    #330.0; DATA = 8'h43;
    #320.0; DATA = 8'h5F;
    #10.0; DATA = 8'hFF;
    #80.0; DATA = 8'h07;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h1E;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'hC2;
    #320.0; DATA = 8'hFF;
    #200.0; DATA = 8'h9E;
    #10.0; DATA = 8'h1E;
    #380.0; DATA = 8'hDE;
    #20.0; DATA = 8'hFA;
    #10.0; DATA = 8'hE2;
    #370.0; DATA = 8'h41;
    #320.0; DATA = 8'hE2;
    #80.0; DATA = 8'h22;
    #10.0; DATA = 8'h26;
    #320.0; DATA = 8'hE2;
    #10.0; DATA = 8'hEB;
    #410.0; DATA = 8'hFF;
    #20.0; DATA = 8'hFA;
    #10.0; DATA = 8'hFF;
    #780.0; DATA = 8'h75;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hF8;
    #330.0; DATA = 8'hFF;
    #320.0; DATA = 8'hC7;
    #10.0; DATA = 8'h43;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'h07;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h1E;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hC2;
    #330.0; DATA = 8'hFF;
    #190.0; DATA = 8'hFE;
    #10.0; DATA = 8'h1E;
    #390.0; DATA = 8'hDE;
    #20.0; DATA = 8'hF2;
    #10.0; DATA = 8'hE2;
    #360.0; DATA = 8'h41;
    #330.0; DATA = 8'hE2;
    #80.0; DATA = 8'h22;
    #10.0; DATA = 8'h26;
    #320.0; DATA = 8'hE2;
    #10.0; DATA = 8'hEF;
    #410.0; DATA = 8'hFF;
    #10.0; DATA = 8'hFE;
    #20.0; DATA = 8'hFF;
    #780.0; DATA = 8'h75;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'hF8;
    #320.0; DATA = 8'hFF;
    #330.0; DATA = 8'h43;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h07;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h1E;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hC2;
    #330.0; DATA = 8'hFF;
    #190.0; DATA = 8'hDE;
    #10.0; DATA = 8'h1E;
    #390.0; DATA = 8'hDE;
    #10.0; DATA = 8'hFA;
    #10.0; DATA = 8'hE2;
    #370.0; DATA = 8'h41;
    #320.0; DATA = 8'h42;
    #10.0; DATA = 8'hE2;
    #80.0; DATA = 8'h26;
    #320.0; DATA = 8'hE2;
    #10.0; DATA = 8'hE3;
    #10.0; DATA = 8'hEB;
    #400.0; DATA = 8'hEF;
    #10.0; DATA = 8'hFF;
    #10.0; DATA = 8'hFA;
    #10.0; DATA = 8'hFF;
    #780.0; DATA = 8'h75;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hF8;
    #330.0; DATA = 8'hFF;
    #330.0; DATA = 8'h43;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h07;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h1E;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'hC2;
    #320.0; DATA = 8'hFF;
    #200.0; DATA = 8'h9E;
    #10.0; DATA = 8'h1E;
    #380.0; DATA = 8'hDE;
    #20.0; DATA = 8'hFA;
    #10.0; DATA = 8'hE2;
    #360.0; DATA = 8'hE0;
    #10.0; DATA = 8'h41;
    #320.0; DATA = 8'hE2;
    #80.0; DATA = 8'h22;
    #10.0; DATA = 8'h26;
    #320.0; DATA = 8'hE2;
    #10.0; DATA = 8'hEB;
    #410.0; DATA = 8'hFF;
    #20.0; DATA = 8'hFA;
    #10.0; DATA = 8'hFF;
    #780.0; DATA = 8'h75;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hF8;
    #330.0; DATA = 8'hFF;
    #320.0; DATA = 8'hF7;
    #10.0; DATA = 8'h43;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'h07;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h1E;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hC2;
    #330.0; DATA = 8'hFF;
    #200.0; DATA = 8'h1E;
    #390.0; DATA = 8'hDE;
    #20.0; DATA = 8'hF2;
    #10.0; DATA = 8'hE2;
    #360.0; DATA = 8'h40;
    #10.0; DATA = 8'h41;
    #320.0; DATA = 8'hE2;
    #80.0; DATA = 8'h22;
    #10.0; DATA = 8'h26;
    #320.0; DATA = 8'hE2;
    #10.0; DATA = 8'hEB;
    #390.0; DATA = 8'hFB;
    #10.0; DATA = 8'hFF;
    #20.0; DATA = 8'hFE;
    #10.0; DATA = 8'hFA;
    #10.0; DATA = 8'hFF;
    #780.0; DATA = 8'h75;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'hF8;
    #320.0; DATA = 8'hFF;
    #330.0; DATA = 8'h43;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h07;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h1E;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hC2;
    #330.0; DATA = 8'hFF;
    #190.0; DATA = 8'hDE;
    #10.0; DATA = 8'h1E;
    #390.0; DATA = 8'hDE;
    #10.0; DATA = 8'hFA;
    #10.0; DATA = 8'hE2;
    #370.0; DATA = 8'h41;
    #330.0; DATA = 8'hE2;
    #80.0; DATA = 8'h26;
    #320.0; DATA = 8'h22;
    #10.0; DATA = 8'hE3;
    #10.0; DATA = 8'hEF;
    #410.0; DATA = 8'hFF;
    #10.0; DATA = 8'hFA;
    #10.0; DATA = 8'hFF;
    #780.0; DATA = 8'h75;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hF8;
    #330.0; DATA = 8'hFF;
    #330.0; DATA = 8'h43;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h07;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h1E;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'hC2;
    #320.0; DATA = 8'hFF;
    #200.0; DATA = 8'h9E;
    #10.0; DATA = 8'h1E;
    #380.0; DATA = 8'hDE;
    #20.0; DATA = 8'hFA;
    #10.0; DATA = 8'hE2;
    #370.0; DATA = 8'h41;
    #320.0; DATA = 8'hE2;
    #80.0; DATA = 8'h22;
    #10.0; DATA = 8'h26;
    #320.0; DATA = 8'hE2;
    #10.0; DATA = 8'hEB;
    #410.0; DATA = 8'hFF;
    #20.0; DATA = 8'hFA;
    #10.0; DATA = 8'hFF;
    #780.0; DATA = 8'h75;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hF8;
    #330.0; DATA = 8'hFF;
    #320.0; DATA = 8'hF7;
    #10.0; DATA = 8'h43;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'h07;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h1E;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hC2;
    #330.0; DATA = 8'hFF;
    #190.0; DATA = 8'hFE;
    #10.0; DATA = 8'h1E;
    #390.0; DATA = 8'hDE;
    #20.0; DATA = 8'hF2;
    #10.0; DATA = 8'hE2;
    #360.0; DATA = 8'h41;
    #330.0; DATA = 8'hE2;
    #460.0; DATA = 8'hEF;
    #10.0; DATA = 8'hAD;
    #400.0; DATA = 8'h81;
    #410.0; DATA = 8'h02;
    #410.0; DATA = 8'h08;
    #410.0; DATA = 8'hCE;
    #410.0; DATA = 8'h66;
    #410.0; DATA = 8'hE2;
    #410.0; DATA = 8'h1E;
    #410.0; DATA = 8'h08;
    #410.0; DATA = 8'hFF;
    #820.0; DATA = 8'hE0;
    #430.0; DATA = 8'h81;
    #330.0; DATA = 8'hE0;
    #90.0; DATA = 8'hF5;
    #320.0; DATA = 8'hE0;
    #10.0; DATA = 8'hFF;
    #70.0; DATA = 8'h12;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hC4;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h2C;
    #320.0; DATA = 8'h2F;
    #10.0; DATA = 8'hFF;
    #350.0; DATA = 8'hFB;
    #10.0; DATA = 8'hE1;
    #10.0; DATA = 8'h01;
    #360.0; DATA = 8'h00;
    #10.0; DATA = 8'h24;
    #320.0; DATA = 8'h01;
    #80.0; DATA = 8'h00;
    #10.0; DATA = 8'hFE;
    #320.0; DATA = 8'h01;
    #10.0; DATA = 8'hFF;
    #150.0; DATA = 8'h3A;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h07;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h78;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h00;
    #330.0; DATA = 8'hFF;
    #220.0; DATA = 8'h00;
    #680.0; DATA = 8'h11;
    #320.0; DATA = 8'h00;
    #20.0; DATA = 8'h02;
    #70.0; DATA = 8'h01;
    #320.0; DATA = 8'h02;
    #10.0; DATA = 8'h23;
    #10.0; DATA = 8'hEF;
    #10.0; DATA = 8'hFF;
    #140.0; DATA = 8'h12;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h07;
    #320.0; DATA = 8'h0F;
    #10.0; DATA = 8'hFF;
    #80.0; DATA = 8'h5F;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h84;
    #320.0; DATA = 8'h9F;
    #10.0; DATA = 8'hFF;
    #570.0; DATA = 8'h24;
    #320.0; DATA = 8'h3F;
    #10.0; DATA = 8'hFF;
    #80.0; DATA = 8'h0F;
    #320.0; DATA = 8'hFF;
    #170.0; DATA = 8'h73;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h01;
    #80.0; DATA = 8'hFF;
    #160.0; DATA = 8'h81;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h3B;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hC4;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h34;
    #330.0; DATA = 8'hFF;
    #380.0; DATA = 8'h00;
    #440.0; DATA = 8'h12;
    #320.0; DATA = 8'h00;
    #10.0; DATA = 8'h01;
    #10.0; DATA = 8'h63;
    #70.0; DATA = 8'hC4;
    #320.0; DATA = 8'h63;
    #10.0; DATA = 8'hFF;
    #70.0; DATA = 8'hBF;
    #10.0; DATA = 8'h08;
    #320.0; DATA = 8'hFF;
    #350.0; DATA = 8'hFB;
    #20.0; DATA = 8'hC1;
    #10.0; DATA = 8'h01;
    #360.0; DATA = 8'h41;
    #10.0; DATA = 8'h73;
    #310.0; DATA = 8'h71;
    #10.0; DATA = 8'h01;
    #80.0; DATA = 8'h0B;
    #10.0; DATA = 8'h3B;
    #70.0; DATA = 8'h01;
    #10.0; DATA = 8'hE3;
    #150.0; DATA = 8'h22;
    #10.0; DATA = 8'h12;
    #320.0; DATA = 8'hE3;
    #10.0; DATA = 8'hFF;
    #80.0; DATA = 8'hC4;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'h27;
    #10.0; DATA = 8'h24;
    #320.0; DATA = 8'hFF;
    #350.0; DATA = 8'hD9;
    #10.0; DATA = 8'h18;
    #10.0; DATA = 8'h00;
    #370.0; DATA = 8'h3A;
    #320.0; DATA = 8'h00;
    #20.0; DATA = 8'h01;
    #70.0; DATA = 8'hC4;
    #320.0; DATA = 8'h01;
    #10.0; DATA = 8'hFF;
    #80.0; DATA = 8'h25;
    #320.0; DATA = 8'hFF;
    #390.0; DATA = 8'h00;
    #440.0; DATA = 8'h12;
    #320.0; DATA = 8'h00;
    #90.0; DATA = 8'hC4;
    #320.0; DATA = 8'h00;
    #10.0; DATA = 8'hEF;
    #10.0; DATA = 8'hFF;
    #60.0; DATA = 8'h23;
    #330.0; DATA = 8'hFF;
    #350.0; DATA = 8'hD8;
    #10.0; DATA = 8'h18;
    #10.0; DATA = 8'h00;
    #370.0; DATA = 8'h3A;
    #320.0; DATA = 8'h00;
    #90.0; DATA = 8'hC4;
    #320.0; DATA = 8'h00;
    #10.0; DATA = 8'hE7;
    #10.0; DATA = 8'hFF;
    #60.0; DATA = 8'h24;
    #330.0; DATA = 8'hFF;
    #390.0; DATA = 8'h00;
    #430.0; DATA = 8'h12;
    #330.0; DATA = 8'h00;
    #80.0; DATA = 8'h07;
    #320.0; DATA = 8'h00;
    #10.0; DATA = 8'hEB;
    #10.0; DATA = 8'hFF;
    #70.0; DATA = 8'h5F;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h81;
    #320.0; DATA = 8'h9F;
    #10.0; DATA = 8'hFF;
    #570.0; DATA = 8'h83;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h24;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h40;
    #320.0; DATA = 8'hFF;
    #170.0; DATA = 8'h93;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h93;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h93;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'h97;
    #10.0; DATA = 8'h93;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'h97;
    #10.0; DATA = 8'h93;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'h93;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h3A;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hC4;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h23;
    #330.0; DATA = 8'hFF;
    #380.0; DATA = 8'h00;
    #440.0; DATA = 8'h12;
    #320.0; DATA = 8'h00;
    #90.0; DATA = 8'h07;
    #320.0; DATA = 8'h00;
    #10.0; DATA = 8'hFF;
    #70.0; DATA = 8'h5F;
    #330.0; DATA = 8'hFF;
    #90.0; DATA = 8'h82;
    #320.0; DATA = 8'hFF;
    #580.0; DATA = 8'h83;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h24;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h40;
    #320.0; DATA = 8'hFF;
    #170.0; DATA = 8'h93;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h93;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'h97;
    #10.0; DATA = 8'h93;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'h93;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h93;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h32;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hC4;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h23;
    #330.0; DATA = 8'hFF;
    #350.0; DATA = 8'hF8;
    #10.0; DATA = 8'h18;
    #10.0; DATA = 8'h00;
    #450.0; DATA = 8'h3A;
    #320.0; DATA = 8'h00;
    #10.0; DATA = 8'h63;
    #10.0; DATA = 8'hE3;
    #60.0; DATA = 8'hC0;
    #10.0; DATA = 8'hC4;
    #320.0; DATA = 8'hE3;
    #10.0; DATA = 8'hFF;
    #70.0; DATA = 8'h23;
    #330.0; DATA = 8'hFF;
    #390.0; DATA = 8'h00;
    #430.0; DATA = 8'h12;
    #330.0; DATA = 8'h00;
    #80.0; DATA = 8'h07;
    #330.0; DATA = 8'h20;
    #10.0; DATA = 8'hF7;
    #10.0; DATA = 8'hFF;
    #60.0; DATA = 8'h5F;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h80;
    #320.0; DATA = 8'h87;
    #10.0; DATA = 8'hFF;
    #570.0; DATA = 8'h83;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h24;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h10;
    #320.0; DATA = 8'hFF;
    #170.0; DATA = 8'h32;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'hC4;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h23;
    #320.0; DATA = 8'hFF;
    #360.0; DATA = 8'hD8;
    #10.0; DATA = 8'h00;
    #460.0; DATA = 8'h3A;
    #320.0; DATA = 8'h00;
    #10.0; DATA = 8'h63;
    #10.0; DATA = 8'hE3;
    #60.0; DATA = 8'hC0;
    #10.0; DATA = 8'hC4;
    #320.0; DATA = 8'hE3;
    #10.0; DATA = 8'hFF;
    #70.0; DATA = 8'h23;
    #330.0; DATA = 8'hFF;
    #380.0; DATA = 8'h80;
    #10.0; DATA = 8'h00;
    #430.0; DATA = 8'h92;
    #320.0; DATA = 8'h00;
    #10.0; DATA = 8'h01;
    #10.0; DATA = 8'h21;
    #10.0; DATA = 8'h61;
    #60.0; DATA = 8'hC4;
    #320.0; DATA = 8'h61;
    #10.0; DATA = 8'hFF;
    #80.0; DATA = 8'h1A;
    #320.0; DATA = 8'hFF;
    #360.0; DATA = 8'hFB;
    #10.0; DATA = 8'hE0;
    #10.0; DATA = 8'h00;
    #360.0; DATA = 8'h60;
    #10.0; DATA = 8'h73;
    #320.0; DATA = 8'h00;
    #10.0; DATA = 8'h40;
    #70.0; DATA = 8'h08;
    #10.0; DATA = 8'h18;
    #320.0; DATA = 8'h40;
    #10.0; DATA = 8'hEB;
    #10.0; DATA = 8'hFF;
    #310.0; DATA = 8'h92;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'hC4;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'h3F;
    #10.0; DATA = 8'h19;
    #320.0; DATA = 8'hFF;
    #350.0; DATA = 8'hFB;
    #20.0; DATA = 8'h00;
    #370.0; DATA = 8'h73;
    #320.0; DATA = 8'h00;
    #20.0; DATA = 8'h20;
    #70.0; DATA = 8'h14;
    #320.0; DATA = 8'h20;
    #10.0; DATA = 8'hEB;
    #10.0; DATA = 8'hEF;
    #10.0; DATA = 8'hFF;
    #300.0; DATA = 8'h92;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hC4;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h1F;
    #330.0; DATA = 8'hFF;
    #350.0; DATA = 8'hFB;
    #10.0; DATA = 8'hFA;
    #10.0; DATA = 8'h00;
    #370.0; DATA = 8'h73;
    #320.0; DATA = 8'h00;
    #10.0; DATA = 8'h20;
    #70.0; DATA = 8'h00;
    #10.0; DATA = 8'h18;
    #320.0; DATA = 8'h20;
    #10.0; DATA = 8'hEB;
    #10.0; DATA = 8'hFF;
    #310.0; DATA = 8'h92;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hC4;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h1E;
    #320.0; DATA = 8'hFF;
    #360.0; DATA = 8'hFB;
    #10.0; DATA = 8'hE0;
    #10.0; DATA = 8'h00;
    #360.0; DATA = 8'h60;
    #10.0; DATA = 8'h73;
    #320.0; DATA = 8'h00;
    #10.0; DATA = 8'h22;
    #70.0; DATA = 8'h00;
    #10.0; DATA = 8'h14;
    #320.0; DATA = 8'h22;
    #10.0; DATA = 8'hFF;
    #320.0; DATA = 8'h13;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'hEF;
    #10.0; DATA = 8'hC4;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'h23;
    #330.0; DATA = 8'hFF;
    #350.0; DATA = 8'hD8;
    #10.0; DATA = 8'h98;
    #10.0; DATA = 8'h00;
    #370.0; DATA = 8'h33;
    #320.0; DATA = 8'h00;
    #90.0; DATA = 8'hC4;
    #320.0; DATA = 8'h00;
    #10.0; DATA = 8'h2B;
    #10.0; DATA = 8'hE3;
    #10.0; DATA = 8'hFF;
    #60.0; DATA = 8'h24;
    #320.0; DATA = 8'hFF;
    #360.0; DATA = 8'hD8;
    #10.0; DATA = 8'h00;
    #460.0; DATA = 8'h84;
    #320.0; DATA = 8'h00;
    #10.0; DATA = 8'h23;
    #80.0; DATA = 8'h27;
    #320.0; DATA = 8'h23;
    #10.0; DATA = 8'hFF;
    #70.0; DATA = 8'hC4;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h25;
    #330.0; DATA = 8'hFF;
    #350.0; DATA = 8'hD8;
    #10.0; DATA = 8'h18;
    #10.0; DATA = 8'h00;
    #450.0; DATA = 8'h25;
    #320.0; DATA = 8'h00;
    #10.0; DATA = 8'h63;
    #70.0; DATA = 8'h03;
    #10.0; DATA = 8'h13;
    #320.0; DATA = 8'h63;
    #10.0; DATA = 8'hFF;
    #160.0; DATA = 8'h73;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h7A;
    #320.0; DATA = 8'hFF;
    #330.0; DATA = 8'h12;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hC4;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h34;
    #330.0; DATA = 8'hFF;
    #350.0; DATA = 8'hD8;
    #10.0; DATA = 8'h18;
    #10.0; DATA = 8'h00;
    #370.0; DATA = 8'h73;
    #320.0; DATA = 8'h00;
    #10.0; DATA = 8'h22;
    #70.0; DATA = 8'h00;
    #10.0; DATA = 8'h05;
    #320.0; DATA = 8'h22;
    #10.0; DATA = 8'hEF;
    #10.0; DATA = 8'hFF;
    #310.0; DATA = 8'h43;
    #320.0; DATA = 8'h4F;
    #10.0; DATA = 8'hFF;
    #80.0; DATA = 8'h07;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h1E;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h82;
    #320.0; DATA = 8'hFF;
    #190.0; DATA = 8'hD8;
    #10.0; DATA = 8'h1C;
    #10.0; DATA = 8'h1E;
    #380.0; DATA = 8'hDE;
    #20.0; DATA = 8'hBE;
    #10.0; DATA = 8'hAE;
    #370.0; DATA = 8'h4D;
    #320.0; DATA = 8'hAE;
    #80.0; DATA = 8'h06;
    #10.0; DATA = 8'h07;
    #320.0; DATA = 8'hAE;
    #10.0; DATA = 8'hEF;
    #70.0; DATA = 8'h3F;
    #10.0; DATA = 8'h1E;
    #320.0; DATA = 8'hEF;
    #10.0; DATA = 8'hFF;
    #70.0; DATA = 8'h81;
    #10.0; DATA = 8'h80;
    #320.0; DATA = 8'hFF;
    #190.0; DATA = 8'hFC;
    #10.0; DATA = 8'h1E;
    #390.0; DATA = 8'hDE;
    #20.0; DATA = 8'hBE;
    #10.0; DATA = 8'hAE;
    #360.0; DATA = 8'h73;
    #330.0; DATA = 8'hAE;
    #10.0; DATA = 8'hAF;
    #70.0; DATA = 8'h02;
    #10.0; DATA = 8'h12;
    #320.0; DATA = 8'hAF;
    #10.0; DATA = 8'hEF;
    #310.0; DATA = 8'hFF;
    #10.0; DATA = 8'h12;
    #320.0; DATA = 8'hEF;
    #10.0; DATA = 8'hFF;
    #80.0; DATA = 8'hC4;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h01;
    #320.0; DATA = 8'hFF;
    #350.0; DATA = 8'hFE;
    #10.0; DATA = 8'hD8;
    #10.0; DATA = 8'h00;
    #370.0; DATA = 8'h73;
    #330.0; DATA = 8'h00;
    #10.0; DATA = 8'h63;
    #70.0; DATA = 8'h1A;
    #320.0; DATA = 8'h43;
    #10.0; DATA = 8'h63;
    #10.0; DATA = 8'hFF;
    #310.0; DATA = 8'h13;
    #10.0; DATA = 8'h12;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'h07;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h5F;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h88;
    #330.0; DATA = 8'hFF;
    #570.0; DATA = 8'h8B;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hC4;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h06;
    #330.0; DATA = 8'hFF;
    #350.0; DATA = 8'hD8;
    #10.0; DATA = 8'hDC;
    #10.0; DATA = 8'h94;
    #340.0; DATA = 8'h95;
    #430.0; DATA = 8'h10;
    #330.0; DATA = 8'h95;
    #80.0; DATA = 8'h81;
    #330.0; DATA = 8'h95;
    #10.0; DATA = 8'hF7;
    #10.0; DATA = 8'hFF;
    #140.0; DATA = 8'h3E;
    #10.0; DATA = 8'h3A;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'hC7;
    #10.0; DATA = 8'hC4;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'h3F;
    #10.0; DATA = 8'h01;
    #320.0; DATA = 8'hFF;
    #390.0; DATA = 8'h81;
    #430.0; DATA = 8'h41;
    #330.0; DATA = 8'h81;
    #80.0; DATA = 8'hC4;
    #320.0; DATA = 8'h81;
    #10.0; DATA = 8'h83;
    #10.0; DATA = 8'hFF;
    #70.0; DATA = 8'h3A;
    #330.0; DATA = 8'hFF;
    #350.0; DATA = 8'hFB;
    #10.0; DATA = 8'hF0;
    #10.0; DATA = 8'h00;
    #380.0; DATA = 8'hFB;
    #20.0; DATA = 8'hE8;
    #370.0; DATA = 8'h54;
    #330.0; DATA = 8'hE8;
    #80.0; DATA = 8'h00;
    #330.0; DATA = 8'hE8;
    #10.0; DATA = 8'hEB;
    #150.0; DATA = 8'h06;
    #330.0; DATA = 8'hEB;
    #10.0; DATA = 8'hFF;
    #70.0; DATA = 8'h24;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hFD;
    #330.0; DATA = 8'hFF;
    #160.0; DATA = 8'h3E;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h10;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h58;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h07;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h5A;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h00;
    #330.0; DATA = 8'hFF;
    #220.0; DATA = 8'hEE;
    #490.0; DATA = 8'h00;
    #680.0; DATA = 8'h41;
    #320.0; DATA = 8'h00;
    #20.0; DATA = 8'h02;
    #70.0; DATA = 8'hC4;
    #320.0; DATA = 8'h02;
    #10.0; DATA = 8'h0B;
    #10.0; DATA = 8'hFF;
    #70.0; DATA = 8'h3C;
    #320.0; DATA = 8'hFF;
    #360.0; DATA = 8'hFB;
    #10.0; DATA = 8'hE1;
    #10.0; DATA = 8'h01;
    #380.0; DATA = 8'hFB;
    #20.0; DATA = 8'hD0;
    #370.0; DATA = 8'h54;
    #330.0; DATA = 8'hD0;
    #80.0; DATA = 8'h00;
    #330.0; DATA = 8'hD0;
    #10.0; DATA = 8'hF3;
    #150.0; DATA = 8'h06;
    #330.0; DATA = 8'hF3;
    #10.0; DATA = 8'hFF;
    #70.0; DATA = 8'h24;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hFD;
    #330.0; DATA = 8'hFF;
    #160.0; DATA = 8'h3E;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h10;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h58;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h07;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h7A;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h00;
    #330.0; DATA = 8'hFF;
    #220.0; DATA = 8'hD6;
    #730.0; DATA = 8'h01;
    #690.0; DATA = 8'h41;
    #320.0; DATA = 8'h01;
    #80.0; DATA = 8'h00;
    #10.0; DATA = 8'hC4;
    #320.0; DATA = 8'h01;
    #10.0; DATA = 8'hFF;
    #70.0; DATA = 8'h3E;
    #330.0; DATA = 8'hFF;
    #350.0; DATA = 8'hFB;
    #20.0; DATA = 8'h00;
    #380.0; DATA = 8'hFB;
    #20.0; DATA = 8'hFF;
    #10.0; DATA = 8'h00;
    #370.0; DATA = 8'h3A;
    #320.0; DATA = 8'h00;
    #90.0; DATA = 8'h07;
    #320.0; DATA = 8'h00;
    #10.0; DATA = 8'hE7;
    #10.0; DATA = 8'hFF;
    #60.0; DATA = 8'h58;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h0C;
    #330.0; DATA = 8'hFF;
    #220.0; DATA = 8'h00;
    #520.0; DATA = 8'h3B;
    #320.0; DATA = 8'h00;
    #20.0; DATA = 8'h63;
    #70.0; DATA = 8'h07;
    #320.0; DATA = 8'h63;
    #10.0; DATA = 8'h6B;
    #10.0; DATA = 8'hFF;
    #70.0; DATA = 8'h78;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h0C;
    #320.0; DATA = 8'hFF;
    #230.0; DATA = 8'h00;
    #510.0; DATA = 8'h12;
    #330.0; DATA = 8'h00;
    #10.0; DATA = 8'h02;
    #70.0; DATA = 8'h00;
    #10.0; DATA = 8'hC4;
    #320.0; DATA = 8'h02;
    #10.0; DATA = 8'hFF;
    #70.0; DATA = 8'h08;
    #330.0; DATA = 8'hFF;
    #350.0; DATA = 8'hFB;
    #20.0; DATA = 8'h01;
    #360.0; DATA = 8'h00;
    #10.0; DATA = 8'h34;
    #320.0; DATA = 8'h01;
    #420.0; DATA = 8'hE3;
    #10.0; DATA = 8'hEF;
    #60.0; DATA = 8'h63;
    #330.0; DATA = 8'hEF;
    #10.0; DATA = 8'hFF;
    #70.0; DATA = 8'h3E;
    #80.0; DATA = 8'hFF;
    #170.0; DATA = 8'h12;
    #320.0; DATA = 8'h13;
    #10.0; DATA = 8'hFF;
    #80.0; DATA = 8'hC4;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h09;
    #320.0; DATA = 8'hFF;
    #350.0; DATA = 8'hFB;
    #20.0; DATA = 8'h83;
    #10.0; DATA = 8'h03;
    #360.0; DATA = 8'h34;
    #330.0; DATA = 8'h03;
    #410.0; DATA = 8'h23;
    #10.0; DATA = 8'hE3;
    #70.0; DATA = 8'h63;
    #320.0; DATA = 8'hE3;
    #10.0; DATA = 8'hFF;
    #80.0; DATA = 8'h37;
    #80.0; DATA = 8'hFF;
    #160.0; DATA = 8'h12;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hC4;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h0A;
    #330.0; DATA = 8'hFF;
    #350.0; DATA = 8'hFB;
    #20.0; DATA = 8'h02;
    #370.0; DATA = 8'h34;
    #320.0; DATA = 8'h02;
    #420.0; DATA = 8'hE3;
    #20.0; DATA = 8'hEB;
    #50.0; DATA = 8'h63;
    #330.0; DATA = 8'hEB;
    #10.0; DATA = 8'hFF;
    #80.0; DATA = 8'h30;
    #80.0; DATA = 8'hFF;
    #160.0; DATA = 8'h38;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h83;
    #330.0; DATA = 8'hFF;
    #160.0; DATA = 8'h8E;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h07;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h09;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h27;
    #330.0; DATA = 8'hFF;
    #180.0; DATA = 8'hFA;
    #10.0; DATA = 8'hD8;
    #10.0; DATA = 8'h26;
    #340.0; DATA = 8'h25;
    #440.0; DATA = 8'h63;
    #320.0; DATA = 8'h25;
    #90.0; DATA = 8'h03;
    #320.0; DATA = 8'h25;
    #20.0; DATA = 8'hEF;
    #10.0; DATA = 8'hFF;
    #300.0; DATA = 8'h41;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hC4;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h26;
    #330.0; DATA = 8'hFF;
    #350.0; DATA = 8'hFD;
    #10.0; DATA = 8'h18;
    #10.0; DATA = 8'h02;
    #380.0; DATA = 8'hDA;
    #20.0; DATA = 8'h1A;
    #10.0; DATA = 8'h02;
    #370.0; DATA = 8'h58;
    #320.0; DATA = 8'h02;
    #80.0; DATA = 8'h00;
    #10.0; DATA = 8'hC4;
    #320.0; DATA = 8'h02;
    #10.0; DATA = 8'hFB;
    #10.0; DATA = 8'hFF;
    #60.0; DATA = 8'h27;
    #330.0; DATA = 8'hFF;
    #390.0; DATA = 8'h02;
    #840.0; DATA = 8'h12;
    #330.0; DATA = 8'h02;
    #80.0; DATA = 8'h07;
    #320.0; DATA = 8'h02;
    #10.0; DATA = 8'h63;
    #10.0; DATA = 8'hFF;
    #70.0; DATA = 8'h09;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h26;
    #320.0; DATA = 8'h3F;
    #10.0; DATA = 8'hFF;
    #180.0; DATA = 8'hFA;
    #10.0; DATA = 8'hDA;
    #10.0; DATA = 8'h02;
    #370.0; DATA = 8'h3A;
    #330.0; DATA = 8'h02;
    #80.0; DATA = 8'hC4;
    #320.0; DATA = 8'h02;
    #10.0; DATA = 8'h03;
    #10.0; DATA = 8'hFB;
    #10.0; DATA = 8'hFF;
    #60.0; DATA = 8'h26;
    #320.0; DATA = 8'h3F;
    #10.0; DATA = 8'hFF;
    #380.0; DATA = 8'h02;
    #440.0; DATA = 8'h8E;
    #320.0; DATA = 8'h02;
    #10.0; DATA = 8'h63;
    #70.0; DATA = 8'h03;
    #10.0; DATA = 8'h07;
    #320.0; DATA = 8'h63;
    #10.0; DATA = 8'hFF;
    #70.0; DATA = 8'h09;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h29;
    #330.0; DATA = 8'hFF;
    #190.0; DATA = 8'hFB;
    #10.0; DATA = 8'hEB;
    #10.0; DATA = 8'h6B;
    #340.0; DATA = 8'h6A;
    #430.0; DATA = 8'h62;
    #10.0; DATA = 8'h63;
    #320.0; DATA = 8'h6A;
    #80.0; DATA = 8'h03;
    #330.0; DATA = 8'h6A;
    #10.0; DATA = 8'hFF;
    #320.0; DATA = 8'h41;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'hC4;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h29;
    #330.0; DATA = 8'hFF;
    #350.0; DATA = 8'hFB;
    #10.0; DATA = 8'hFA;
    #10.0; DATA = 8'h00;
    #380.0; DATA = 8'hFB;
    #30.0; DATA = 8'h00;
    #370.0; DATA = 8'h58;
    #320.0; DATA = 8'h00;
    #90.0; DATA = 8'hC4;
    #320.0; DATA = 8'h00;
    #10.0; DATA = 8'hEB;
    #10.0; DATA = 8'hFB;
    #10.0; DATA = 8'hFF;
    #50.0; DATA = 8'h2A;
    #330.0; DATA = 8'hFF;
    #390.0; DATA = 8'h00;
    #840.0; DATA = 8'h12;
    #330.0; DATA = 8'h00;
    #80.0; DATA = 8'h07;
    #330.0; DATA = 8'h20;
    #10.0; DATA = 8'hF7;
    #10.0; DATA = 8'hFF;
    #60.0; DATA = 8'h09;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h28;
    #330.0; DATA = 8'hFF;
    #180.0; DATA = 8'hFB;
    #20.0; DATA = 8'h00;
    #370.0; DATA = 8'h3A;
    #320.0; DATA = 8'h00;
    #90.0; DATA = 8'hC4;
    #320.0; DATA = 8'h80;
    #10.0; DATA = 8'h01;
    #10.0; DATA = 8'hE3;
    #10.0; DATA = 8'hFF;
    #60.0; DATA = 8'h29;
    #320.0; DATA = 8'hFF;
    #390.0; DATA = 8'h00;
    #440.0; DATA = 8'h60;
    #320.0; DATA = 8'h00;
    #90.0; DATA = 8'h1C;
    #320.0; DATA = 8'h00;
    #10.0; DATA = 8'hFD;
    #10.0; DATA = 8'hFF;
    #310.0; DATA = 8'h12;
    #320.0; DATA = 8'h1B;
    #10.0; DATA = 8'hFF;
    #80.0; DATA = 8'hC4;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h2C;
    #320.0; DATA = 8'hFF;
    #350.0; DATA = 8'hFB;
    #20.0; DATA = 8'hE1;
    #10.0; DATA = 8'h01;
    #360.0; DATA = 8'h20;
    #10.0; DATA = 8'h3A;
    #320.0; DATA = 8'h01;
    #10.0; DATA = 8'h21;
    #70.0; DATA = 8'h05;
    #10.0; DATA = 8'h07;
    #320.0; DATA = 8'h21;
    #10.0; DATA = 8'hFF;
    #70.0; DATA = 8'h78;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h00;
    #330.0; DATA = 8'hFF;
    #220.0; DATA = 8'h01;
    #510.0; DATA = 8'h00;
    #10.0; DATA = 8'h12;
    #320.0; DATA = 8'h01;
    #10.0; DATA = 8'h21;
    #70.0; DATA = 8'h00;
    #10.0; DATA = 8'hC4;
    #320.0; DATA = 8'h21;
    #10.0; DATA = 8'hFF;
    #70.0; DATA = 8'h08;
    #330.0; DATA = 8'hFF;
    #350.0; DATA = 8'hFB;
    #20.0; DATA = 8'h01;
    #360.0; DATA = 8'h00;
    #10.0; DATA = 8'h9C;
    #320.0; DATA = 8'h01;
    #10.0; DATA = 8'h21;
    #70.0; DATA = 8'h00;
    #10.0; DATA = 8'h42;
    #320.0; DATA = 8'h21;
    #10.0; DATA = 8'hFF;
    #70.0; DATA = 8'hE4;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h4F;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hA9;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hA8;
    #330.0; DATA = 8'hFF;
    #490.0; DATA = 8'h8A;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hA7;
    #320.0; DATA = 8'hBF;
    #10.0; DATA = 8'hFF;
    #220.0; DATA = 8'h29;
    #400.0; DATA = 8'hAD;
    #10.0; DATA = 8'h84;
    #430.0; DATA = 8'h13;
    #320.0; DATA = 8'h17;
    #10.0; DATA = 8'h84;
    #10.0; DATA = 8'hA7;
    #70.0; DATA = 8'hC4;
    #320.0; DATA = 8'h84;
    #10.0; DATA = 8'hA7;
    #10.0; DATA = 8'hFF;
    #70.0; DATA = 8'h02;
    #330.0; DATA = 8'hFF;
    #350.0; DATA = 8'hD8;
    #10.0; DATA = 8'h14;
    #10.0; DATA = 8'h00;
    #370.0; DATA = 8'h7B;
    #320.0; DATA = 8'h00;
    #10.0; DATA = 8'h63;
    #70.0; DATA = 8'h00;
    #330.0; DATA = 8'h63;
    #10.0; DATA = 8'hEF;
    #70.0; DATA = 8'hD8;
    #330.0; DATA = 8'hEF;
    #10.0; DATA = 8'hFF;
    #150.0; DATA = 8'h12;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hC4;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h09;
    #330.0; DATA = 8'hFF;
    #350.0; DATA = 8'hFB;
    #20.0; DATA = 8'h03;
    #360.0; DATA = 8'h02;
    #10.0; DATA = 8'h9C;
    #320.0; DATA = 8'h03;
    #10.0; DATA = 8'h23;
    #10.0; DATA = 8'h63;
    #60.0; DATA = 8'h42;
    #330.0; DATA = 8'h63;
    #10.0; DATA = 8'hE3;
    #70.0; DATA = 8'hE0;
    #10.0; DATA = 8'hE4;
    #320.0; DATA = 8'hE3;
    #10.0; DATA = 8'hFF;
    #70.0; DATA = 8'hE0;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hA8;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hA8;
    #330.0; DATA = 8'hFF;
    #490.0; DATA = 8'h8D;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hD5;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h12;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hC4;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h0A;
    #330.0; DATA = 8'hFF;
    #350.0; DATA = 8'hFB;
    #10.0; DATA = 8'hF3;
    #10.0; DATA = 8'h02;
    #360.0; DATA = 8'h00;
    #10.0; DATA = 8'h9C;
    #320.0; DATA = 8'h02;
    #90.0; DATA = 8'h42;
    #320.0; DATA = 8'h02;
    #10.0; DATA = 8'hE3;
    #10.0; DATA = 8'hEB;
    #60.0; DATA = 8'hE1;
    #10.0; DATA = 8'hE5;
    #320.0; DATA = 8'hEB;
    #10.0; DATA = 8'hFF;
    #70.0; DATA = 8'h02;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hA8;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hA8;
    #330.0; DATA = 8'hFF;
    #490.0; DATA = 8'h8E;
    #320.0; DATA = 8'h8F;
    #10.0; DATA = 8'hFF;
    #80.0; DATA = 8'h69;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h12;
    #320.0; DATA = 8'hDF;
    #10.0; DATA = 8'hFF;
    #80.0; DATA = 8'hC4;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h29;
    #320.0; DATA = 8'hFF;
    #350.0; DATA = 8'hFB;
    #20.0; DATA = 8'hC0;
    #10.0; DATA = 8'h00;
    #360.0; DATA = 8'h28;
    #330.0; DATA = 8'h00;
    #80.0; DATA = 8'h80;
    #320.0; DATA = 8'h00;
    #10.0; DATA = 8'h23;
    #10.0; DATA = 8'hE3;
    #10.0; DATA = 8'hFF;
    #140.0; DATA = 8'h73;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h3A;
    #330.0; DATA = 8'hFF;
    #320.0; DATA = 8'h17;
    #10.0; DATA = 8'h12;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'hC4;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h06;
    #330.0; DATA = 8'hFF;
    #350.0; DATA = 8'hD8;
    #10.0; DATA = 8'hDC;
    #10.0; DATA = 8'h95;
    #370.0; DATA = 8'h28;
    #320.0; DATA = 8'h95;
    #90.0; DATA = 8'h1F;
    #320.0; DATA = 8'h95;
    #10.0; DATA = 8'hF7;
    #10.0; DATA = 8'hFF;
    #150.0; DATA = 8'h73;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h04;
    #80.0; DATA = 8'hFF;
    #160.0; DATA = 8'h24;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h20;
    #330.0; DATA = 8'hFF;
    #160.0; DATA = 8'hAA;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h5F;
    #330.0; DATA = 8'hFF;
    #300.0; DATA = 8'hB5;
    #410.0; DATA = 8'h8E;
    #440.0; DATA = 8'h42;
    #320.0; DATA = 8'h8E;
    #80.0; DATA = 8'h04;
    #10.0; DATA = 8'h44;
    #320.0; DATA = 8'h8E;
    #10.0; DATA = 8'hFF;
    #70.0; DATA = 8'h19;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h46;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hE5;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h08;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h12;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h50;
    #330.0; DATA = 8'hFF;
    #410.0; DATA = 8'hA7;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h73;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h15;
    #80.0; DATA = 8'hFF;
    #160.0; DATA = 8'h34;
    #330.0; DATA = 8'hFF;
    #490.0; DATA = 8'h73;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h16;
    #80.0; DATA = 8'hFF;
    #160.0; DATA = 8'h3A;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h25;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h20;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h00;
    #330.0; DATA = 8'hFF;
    #300.0; DATA = 8'hA7;
    #680.0; DATA = 8'h12;
    #330.0; DATA = 8'hA7;
    #80.0; DATA = 8'h50;
    #330.0; DATA = 8'hA7;
    #10.0; DATA = 8'hFF;
    #400.0; DATA = 8'hB7;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h3A;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h25;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h20;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'hC1;
    #10.0; DATA = 8'h40;
    #320.0; DATA = 8'hFF;
    #300.0; DATA = 8'hB7;
    #520.0; DATA = 8'h82;
    #330.0; DATA = 8'hB7;
    #80.0; DATA = 8'h24;
    #320.0; DATA = 8'h37;
    #10.0; DATA = 8'hF7;
    #80.0; DATA = 8'h40;
    #320.0; DATA = 8'h43;
    #10.0; DATA = 8'hFF;
    #540.0; DATA = 8'h00;
    #600.0; DATA = 8'h82;
    #330.0; DATA = 8'h00;
    #80.0; DATA = 8'h20;
    #330.0; DATA = 8'h02;
    #10.0; DATA = 8'hE3;
    #10.0; DATA = 8'hFF;
    #440.0; DATA = 8'h00;
    #770.0; DATA = 8'h60;
    #320.0; DATA = 8'h00;
    #90.0; DATA = 8'hE7;
    #320.0; DATA = 8'h00;
    #10.0; DATA = 8'hE7;
    #10.0; DATA = 8'hFF;
    #310.0; DATA = 8'h12;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h50;
    #320.0; DATA = 8'hFF;
    #410.0; DATA = 8'h01;
    #10.0; DATA = 8'h00;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'h73;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h15;
    #330.0; DATA = 8'hFF;
    #330.0; DATA = 8'h08;
    #320.0; DATA = 8'h0B;
    #10.0; DATA = 8'hFF;
    #80.0; DATA = 8'h24;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h01;
    #320.0; DATA = 8'hFF;
    #740.0; DATA = 8'h60;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hE2;
    #330.0; DATA = 8'hFF;
    #320.0; DATA = 8'h1F;
    #10.0; DATA = 8'h12;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'h50;
    #330.0; DATA = 8'hFF;
    #410.0; DATA = 8'hED;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h73;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h15;
    #80.0; DATA = 8'hFF;
    #160.0; DATA = 8'h34;
    #330.0; DATA = 8'hFF;
    #490.0; DATA = 8'h73;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h16;
    #80.0; DATA = 8'hFF;
    #170.0; DATA = 8'h3A;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h25;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h20;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h00;
    #320.0; DATA = 8'hFF;
    #300.0; DATA = 8'hED;
    #600.0; DATA = 8'h12;
    #330.0; DATA = 8'hED;
    #10.0; DATA = 8'hEF;
    #70.0; DATA = 8'h50;
    #330.0; DATA = 8'hEF;
    #10.0; DATA = 8'hFF;
    #400.0; DATA = 8'hFD;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h3A;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h25;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h20;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h40;
    #320.0; DATA = 8'hFF;
    #300.0; DATA = 8'hFD;
    #520.0; DATA = 8'h82;
    #330.0; DATA = 8'hFD;
    #80.0; DATA = 8'h24;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h40;
    #330.0; DATA = 8'hFF;
    #540.0; DATA = 8'hBF;
    #10.0; DATA = 8'h00;
    #590.0; DATA = 8'h82;
    #330.0; DATA = 8'h00;
    #80.0; DATA = 8'h20;
    #330.0; DATA = 8'h00;
    #10.0; DATA = 8'hA3;
    #10.0; DATA = 8'hFF;
    #440.0; DATA = 8'h00;
    #770.0; DATA = 8'h60;
    #320.0; DATA = 8'h00;
    #90.0; DATA = 8'hE7;
    #320.0; DATA = 8'h00;
    #10.0; DATA = 8'hE7;
    #10.0; DATA = 8'hFF;
    #310.0; DATA = 8'h12;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h50;
    #330.0; DATA = 8'hFF;
    #400.0; DATA = 8'hAF;
    #10.0; DATA = 8'h00;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'h77;
    #10.0; DATA = 8'h73;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'h15;
    #330.0; DATA = 8'hFF;
    #330.0; DATA = 8'h08;
    #320.0; DATA = 8'h0B;
    #10.0; DATA = 8'hFF;
    #80.0; DATA = 8'h24;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h01;
    #320.0; DATA = 8'hFF;
    #740.0; DATA = 8'h60;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hE2;
    #330.0; DATA = 8'hFF;
    #320.0; DATA = 8'h1F;
    #10.0; DATA = 8'h12;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'h50;
    #330.0; DATA = 8'hFF;
    #410.0; DATA = 8'hEA;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h73;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h15;
    #80.0; DATA = 8'hFF;
    #160.0; DATA = 8'h34;
    #330.0; DATA = 8'hFF;
    #490.0; DATA = 8'h73;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h16;
    #80.0; DATA = 8'hFF;
    #170.0; DATA = 8'h3A;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'h27;
    #10.0; DATA = 8'h25;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h20;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'h00;
    #330.0; DATA = 8'hFF;
    #300.0; DATA = 8'hEA;
    #600.0; DATA = 8'h12;
    #330.0; DATA = 8'hEA;
    #80.0; DATA = 8'h50;
    #330.0; DATA = 8'hEA;
    #10.0; DATA = 8'hFF;
    #400.0; DATA = 8'hFA;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h3A;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h25;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h20;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'hC7;
    #10.0; DATA = 8'h40;
    #320.0; DATA = 8'hFF;
    #300.0; DATA = 8'hFA;
    #520.0; DATA = 8'h82;
    #330.0; DATA = 8'hFA;
    #80.0; DATA = 8'h24;
    #320.0; DATA = 8'h20;
    #10.0; DATA = 8'hFB;
    #10.0; DATA = 8'hFF;
    #70.0; DATA = 8'h40;
    #330.0; DATA = 8'hFF;
    #540.0; DATA = 8'hBF;
    #10.0; DATA = 8'h00;
    #590.0; DATA = 8'h82;
    #330.0; DATA = 8'h00;
    #80.0; DATA = 8'h20;
    #330.0; DATA = 8'h00;
    #10.0; DATA = 8'hA3;
    #10.0; DATA = 8'hFF;
    #440.0; DATA = 8'h00;
    #770.0; DATA = 8'h60;
    #320.0; DATA = 8'h00;
    #90.0; DATA = 8'hE7;
    #320.0; DATA = 8'h00;
    #10.0; DATA = 8'hE7;
    #10.0; DATA = 8'hFF;
    #310.0; DATA = 8'h12;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h50;
    #330.0; DATA = 8'hFF;
    #400.0; DATA = 8'hBF;
    #10.0; DATA = 8'h00;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'hF7;
    #10.0; DATA = 8'h73;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'h15;
    #330.0; DATA = 8'hFF;
    #330.0; DATA = 8'h08;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h24;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h01;
    #320.0; DATA = 8'hFF;
    #740.0; DATA = 8'h60;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'hE2;
    #330.0; DATA = 8'hFF;
    #320.0; DATA = 8'h3F;
    #10.0; DATA = 8'h12;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'h50;
    #330.0; DATA = 8'hFF;
    #410.0; DATA = 8'h88;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h73;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h15;
    #80.0; DATA = 8'hFF;
    #160.0; DATA = 8'h34;
    #330.0; DATA = 8'hFF;
    #490.0; DATA = 8'h73;
    #330.0; DATA = 8'hFF;
    #80.0; DATA = 8'h16;
    #80.0; DATA = 8'hFF;
    #170.0; DATA = 8'h3A;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'hE7;
    #10.0; DATA = 8'h25;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h20;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'h05;
    #10.0; DATA = 8'h00;
    #320.0; DATA = 8'hFF;
    #300.0; DATA = 8'h88;
    #600.0; DATA = 8'h12;
    #330.0; DATA = 8'h88;
    #10.0; DATA = 8'hAB;
    #70.0; DATA = 8'h00;
    #10.0; DATA = 8'h50;
    #320.0; DATA = 8'hAB;
    #10.0; DATA = 8'hFF;
    #400.0; DATA = 8'h98;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h3A;
    #320.0; DATA = 8'hFF;
    #90.0; DATA = 8'h25;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'hFA;
    #10.0; DATA = 8'h20;
    #320.0; DATA = 8'hFF;
    #80.0; DATA = 8'h40;
    #330.0; DATA = 8'hFF;
    #300.0; DATA = 8'h98;
    #520.0; DATA = 8'h82;
    #320.0; DATA = 8'h88;
    #10.0; DATA = 8'h98;
    #80.0; DATA = 8'h24;
    #320.0; DATA = 8'h98;
    #10.0; DATA = 8'h9B;
    #10.0; DATA = 8'hFF;
    #70.0; DATA = 8'h40;
    #320.0; DATA = 8'h41;
    #10.0; DATA = 8'hFF;
    #540.0; DATA = 8'h00;
    #600.0; DATA = 8'h82;
    #330.0; DATA = 8'h00;
    #80.0; DATA = 8'h20;
    #330.0; DATA = 8'h00;
    #10.0; DATA = 8'hA3;
    #10.0; DATA = 8'hFF;
    #440.0; DATA = 8'h00;

end
initial
begin
    RWb = 1'b1;
    #60550.0; RWb = 1'b0;
    #4910.0; RWb = 1'b1;
    #5400.0; RWb = 1'b0;
    #660.0; RWb = 1'b1;
    #6540.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #5980.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #3440.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #7450.0; RWb = 1'b0;
    #400.0; RWb = 1'b1;
    #9010.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #6960.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #36010.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #2460.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #7120.0; RWb = 1'b0;
    #1150.0; RWb = 1'b1;
    #7120.0; RWb = 1'b0;
    #1390.0; RWb = 1'b1;
    #4090.0; RWb = 1'b0;
    #500.0; RWb = 1'b1;
    #1800.0; RWb = 1'b0;
    #490.0; RWb = 1'b1;
    #13100.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #4910.0; RWb = 1'b0;
    #820.0; RWb = 1'b1;
    #3680.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #2130.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #4910.0; RWb = 1'b0;
    #820.0; RWb = 1'b1;
    #3680.0; RWb = 1'b0;
    #410.0; RWb = 1'b1;
    #4750.0; RWb = 1'b0;
    #490.0; RWb = 1'b1;
    #5730.0; RWb = 1'b0;
    #820.0; RWb = 1'b1;
    #23570.0; RWb = 1'b0;
    #820.0; RWb = 1'b1;
    #8020.0; RWb = 1'b0;
    #660.0; RWb = 1'b1;
    #3440.0; RWb = 1'b0;
    #490.0; RWb = 1'b1;
    #1720.0; RWb = 1'b0;
    #570.0; RWb = 1'b1;
    #1230.0; RWb = 1'b0;
    #730.0; RWb = 1'b1;
    #12200.0; RWb = 1'b0;
    #570.0; RWb = 1'b1;
    #3440.0; RWb = 1'b0;
    #490.0; RWb = 1'b1;
    #1720.0; RWb = 1'b0;
    #570.0; RWb = 1'b1;
    #1230.0; RWb = 1'b0;
    #730.0; RWb = 1'b1;
    #12200.0; RWb = 1'b0;
    #570.0; RWb = 1'b1;
    #3440.0; RWb = 1'b0;
    #490.0; RWb = 1'b1;
    #1720.0; RWb = 1'b0;
    #570.0; RWb = 1'b1;
    #1230.0; RWb = 1'b0;
    #730.0; RWb = 1'b1;
    #12200.0; RWb = 1'b0;
    #570.0; RWb = 1'b1;
    #3440.0; RWb = 1'b0;
    #490.0; RWb = 1'b1;
    #1720.0; RWb = 1'b0;
    #570.0; RWb = 1'b1;
    #1230.0; RWb = 1'b0;

end
initial
begin
    AS2 = 1'b0;
    #30.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #170.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #410.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #410.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #170.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #410.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #170.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #410.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #410.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #170.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #420.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #170.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #410.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #410.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #410.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #170.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #410.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #490.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #240.0; AS2 = 1'b0;
    #580.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #170.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #170.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #170.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #80.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #410.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #80.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #410.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #410.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #170.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #170.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #410.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #170.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #170.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #170.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #410.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #170.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #170.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #410.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #170.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #170.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #170.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #410.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #320.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #250.0; AS2 = 1'b0;
    #410.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #570.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #250.0; AS2 = 1'b0;
    #660.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #570.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #250.0; AS2 = 1'b0;
    #400.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #250.0; AS2 = 1'b0;
    #410.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #80.0; AS2 = 1'b1;
    #170.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #80.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #90.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #410.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #170.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #410.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #410.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #420.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #250.0; AS2 = 1'b0;
    #410.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #490.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #250.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #490.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #320.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #490.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #170.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #320.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #170.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #80.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #410.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #80.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #80.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #570.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #410.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #410.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #580.0; AS2 = 1'b0;
    #490.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #490.0; AS2 = 1'b0;
    #650.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #410.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #740.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #320.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #410.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #80.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #80.0; AS2 = 1'b1;
    #170.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #490.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #410.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #410.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #570.0; AS2 = 1'b0;
    #490.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #490.0; AS2 = 1'b0;
    #650.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #420.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #740.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #320.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #410.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #80.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #80.0; AS2 = 1'b1;
    #170.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #490.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #410.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #410.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #580.0; AS2 = 1'b0;
    #490.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #490.0; AS2 = 1'b0;
    #650.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #420.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #740.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #320.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #410.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #80.0; AS2 = 1'b1;
    #160.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #80.0; AS2 = 1'b1;
    #170.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #490.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #410.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #330.0; AS2 = 1'b0;
    #410.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #90.0; AS2 = 1'b0;
    #320.0; AS2 = 1'b1;
    #580.0; AS2 = 1'b0;
    #490.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #80.0; AS2 = 1'b0;
    #330.0; AS2 = 1'b1;
    #490.0; AS2 = 1'b0;

end
initial
begin
    DTAC2 = 1'b0;
    #50.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #620.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #620.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #320.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #540.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #540.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #440.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #460.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #540.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #570.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #330.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #690.0; DTAC2 = 1'b0;
    #90.0; DTAC2 = 1'b1;
    #570.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #330.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #330.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #330.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #540.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #330.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #370.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #620.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #280.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #290.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #700.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #330.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #540.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #320.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #330.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #940.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #330.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #850.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #610.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #330.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #330.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #330.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #940.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #330.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #850.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #620.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #330.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #540.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #320.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #330.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #940.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #330.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #450.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #620.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #330.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #530.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #210.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #540.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #320.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;
    #860.0; DTAC2 = 1'b0;
    #80.0; DTAC2 = 1'b1;
    #330.0; DTAC2 = 1'b0;
    #200.0; DTAC2 = 1'b1;
    #200.0; DTAC2 = 1'b0;
    #210.0; DTAC2 = 1'b1;

end
initial
begin
    VRAMCS2 = 1'b1;
    #71150.0; VRAMCS2 = 1'b0;
    #10.0; VRAMCS2 = 1'b1;
    #88720.0; VRAMCS2 = 1'b0;
    #370.0; VRAMCS2 = 1'b1;
    #290.0; VRAMCS2 = 1'b0;
    #370.0; VRAMCS2 = 1'b1;
    #7490.0; VRAMCS2 = 1'b0;
    #370.0; VRAMCS2 = 1'b1;
    #280.0; VRAMCS2 = 1'b0;
    #380.0; VRAMCS2 = 1'b1;
    #4210.0; VRAMCS2 = 1'b0;
    #370.0; VRAMCS2 = 1'b1;
    #1920.0; VRAMCS2 = 1'b0;
    #370.0; VRAMCS2 = 1'b1;
    #40560.0; VRAMCS2 = 1'b0;
    #10.0; VRAMCS2 = 1'b1;
    #39610.0; VRAMCS2 = 1'b0;
    #370.0; VRAMCS2 = 1'b1;
    #3560.0; VRAMCS2 = 1'b0;
    #370.0; VRAMCS2 = 1'b1;
    #1920.0; VRAMCS2 = 1'b0;
    #370.0; VRAMCS2 = 1'b1;
    #1590.0; VRAMCS2 = 1'b0;
    #380.0; VRAMCS2 = 1'b1;
    #12390.0; VRAMCS2 = 1'b0;
    #370.0; VRAMCS2 = 1'b1;
    #3560.0; VRAMCS2 = 1'b0;
    #370.0; VRAMCS2 = 1'b1;
    #1920.0; VRAMCS2 = 1'b0;
    #370.0; VRAMCS2 = 1'b1;
    #1590.0; VRAMCS2 = 1'b0;
    #380.0; VRAMCS2 = 1'b1;
    #12390.0; VRAMCS2 = 1'b0;
    #370.0; VRAMCS2 = 1'b1;
    #3560.0; VRAMCS2 = 1'b0;
    #370.0; VRAMCS2 = 1'b1;
    #1920.0; VRAMCS2 = 1'b0;
    #370.0; VRAMCS2 = 1'b1;
    #1590.0; VRAMCS2 = 1'b0;
    #380.0; VRAMCS2 = 1'b1;
    #12390.0; VRAMCS2 = 1'b0;
    #370.0; VRAMCS2 = 1'b1;
    #3560.0; VRAMCS2 = 1'b0;
    #370.0; VRAMCS2 = 1'b1;
    #1920.0; VRAMCS2 = 1'b0;
    #370.0; VRAMCS2 = 1'b1;
    #1590.0; VRAMCS2 = 1'b0;

end
initial
begin
    #330000.0; $finish;
end
endmodule